// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.1.0.96
// Netlist written on Sat Sep 27 02:20:49 2014
//
// Verilog Description of module main
//

module main (SCLK, MOSI, MISO, CE1, GSRn, SDA);   // c:/users/yisong/documents/new/mlp/main.vhd(20[8:12])
    input SCLK /* synthesis black_box_pad_pin=1 */ ;   // c:/users/yisong/documents/new/mlp/main.vhd(21[8:12])
    input MOSI /* synthesis black_box_pad_pin=1 */ ;   // c:/users/yisong/documents/new/mlp/main.vhd(22[4:8])
    output MISO /* synthesis black_box_pad_pin=1 */ ;   // c:/users/yisong/documents/new/mlp/main.vhd(23[4:8])
    input CE1;   // c:/users/yisong/documents/new/mlp/main.vhd(24[4:7])
    input GSRn;   // c:/users/yisong/documents/new/mlp/main.vhd(25[4:8])
    input SDA;   // c:/users/yisong/documents/new/mlp/main.vhd(44[4:7])
    
    wire [31:0]inputNumber;   // c:/users/yisong/documents/new/mlp/loadweight.vhd(22[2:13])
    wire CE1_c;   // c:/users/yisong/documents/new/mlp/main.vhd(24[4:7])
    wire SDA_c;   // c:/users/yisong/documents/new/mlp/main.vhd(44[4:7])
    wire GSRnX /* synthesis pullmode="UP" */ ;   // c:/users/yisong/documents/new/mlp/main.vhd(246[8:13])
    wire clock;   // c:/users/yisong/documents/new/mlp/main.vhd(251[8:13])
    wire [7:0]writeout;   // c:/users/yisong/documents/new/mlp/main.vhd(253[8:16])
    wire [7:0]write_data;   // c:/users/yisong/documents/new/mlp/main.vhd(260[8:18])
    wire [7:0]read_data;   // c:/users/yisong/documents/new/mlp/main.vhd(262[8:17])
    wire new_data;   // c:/users/yisong/documents/new/mlp/main.vhd(263[8:16])
    wire [31:0]ramDataIn;   // c:/users/yisong/documents/new/mlp/main.vhd(272[8:17])
    wire weight_done;   // c:/users/yisong/documents/new/mlp/main.vhd(277[8:19])
    wire [11:0]sram_address_A;   // c:/users/yisong/documents/new/mlp/main.vhd(281[8:22])
    wire [31:0]sram_input_A;   // c:/users/yisong/documents/new/mlp/main.vhd(282[8:20])
    wire sram_ready_A;   // c:/users/yisong/documents/new/mlp/main.vhd(285[8:20])
    wire [11:0]sram_address_B;   // c:/users/yisong/documents/new/mlp/main.vhd(288[8:22])
    wire [31:0]sram_output_B;   // c:/users/yisong/documents/new/mlp/main.vhd(290[8:21])
    wire sram_ready_B;   // c:/users/yisong/documents/new/mlp/main.vhd(292[8:20])
    wire float_alu_ready;   // c:/users/yisong/documents/new/mlp/main.vhd(296[8:23])
    wire [31:0]float_alu_b;   // c:/users/yisong/documents/new/mlp/main.vhd(297[21:32])
    wire [31:0]float_alu_c;   // c:/users/yisong/documents/new/mlp/main.vhd(297[34:45])
    wire [2:0]float_alu_mode;   // c:/users/yisong/documents/new/mlp/main.vhd(298[8:22])
    wire [31:0]\mlp_outputs[1] ;   // c:/users/yisong/documents/new/mlp/main.vhd(302[8:19])
    wire [31:0]\mlp_outputs[0] ;   // c:/users/yisong/documents/new/mlp/main.vhd(302[8:19])
    wire mlp_done;   // c:/users/yisong/documents/new/mlp/main.vhd(304[8:16])
    wire output_new;   // c:/users/yisong/documents/new/mlp/main.vhd(312[8:18])
    wire [31:0]count;   // c:/users/yisong/documents/new/mlp/receiver.vhd(20[8:13])
    wire [31:0]i;   // c:/users/yisong/documents/new/mlp/test.vhd(166[8:9])
    wire [3:0]n236;   // mult_2u_2u.v(11[23:24])
    wire mco_131;   // mult_24u_24u.v(944[10:17])
    wire mult_24u_24u_0_pp_11_45;   // mult_24u_24u.v(943[10:33])
    wire mult_24u_24u_0_pp_11_46;   // mult_24u_24u.v(942[10:33])
    wire mfco_11;   // mult_24u_24u.v(941[10:17])
    wire mco_130;   // mult_24u_24u.v(940[10:17])
    wire mult_24u_24u_0_pp_11_43;   // mult_24u_24u.v(939[10:33])
    wire mult_24u_24u_0_pp_11_44;   // mult_24u_24u.v(938[10:33])
    wire mco_129;   // mult_24u_24u.v(937[10:17])
    wire mult_24u_24u_0_pp_11_41;   // mult_24u_24u.v(936[10:33])
    wire mult_24u_24u_0_pp_11_42;   // mult_24u_24u.v(935[10:33])
    wire mco_128;   // mult_24u_24u.v(934[10:17])
    wire mult_24u_24u_0_pp_11_39;   // mult_24u_24u.v(933[10:33])
    wire mult_24u_24u_0_pp_11_40;   // mult_24u_24u.v(932[10:33])
    wire mco_127;   // mult_24u_24u.v(931[10:17])
    wire mult_24u_24u_0_pp_11_37;   // mult_24u_24u.v(930[10:33])
    wire mult_24u_24u_0_pp_11_38;   // mult_24u_24u.v(929[10:33])
    wire mco_126;   // mult_24u_24u.v(928[10:17])
    wire mult_24u_24u_0_pp_11_35;   // mult_24u_24u.v(927[10:33])
    wire mult_24u_24u_0_pp_11_36;   // mult_24u_24u.v(926[10:33])
    wire mco_125;   // mult_24u_24u.v(925[10:17])
    wire mult_24u_24u_0_pp_11_33;   // mult_24u_24u.v(924[10:33])
    wire mult_24u_24u_0_pp_11_34;   // mult_24u_24u.v(923[10:33])
    wire mco_124;   // mult_24u_24u.v(922[10:17])
    wire mult_24u_24u_0_pp_11_31;   // mult_24u_24u.v(921[10:33])
    wire mult_24u_24u_0_pp_11_32;   // mult_24u_24u.v(920[10:33])
    wire mco_123;   // mult_24u_24u.v(919[10:17])
    wire mult_24u_24u_0_pp_11_29;   // mult_24u_24u.v(918[10:33])
    wire mult_24u_24u_0_pp_11_30;   // mult_24u_24u.v(917[10:33])
    wire mco_122;   // mult_24u_24u.v(916[10:17])
    wire mult_24u_24u_0_pp_11_27;   // mult_24u_24u.v(915[10:33])
    wire mult_24u_24u_0_pp_11_28;   // mult_24u_24u.v(914[10:33])
    wire mco_121;   // mult_24u_24u.v(913[10:17])
    wire mult_24u_24u_0_pp_11_25;   // mult_24u_24u.v(912[10:33])
    wire mult_24u_24u_0_pp_11_26;   // mult_24u_24u.v(911[10:33])
    wire mult_24u_24u_0_cin_lr_22;   // mult_24u_24u.v(910[10:34])
    wire mult_24u_24u_0_pp_11_23;   // mult_24u_24u.v(909[10:33])
    wire mult_24u_24u_0_pp_11_24;   // mult_24u_24u.v(908[10:33])
    wire mco_120;   // mult_24u_24u.v(907[10:17])
    wire mult_24u_24u_0_pp_10_43;   // mult_24u_24u.v(906[10:33])
    wire mult_24u_24u_0_pp_10_44;   // mult_24u_24u.v(905[10:33])
    wire mfco_10;   // mult_24u_24u.v(904[10:17])
    wire mco_119;   // mult_24u_24u.v(903[10:17])
    wire mult_24u_24u_0_pp_10_41;   // mult_24u_24u.v(902[10:33])
    wire mult_24u_24u_0_pp_10_42;   // mult_24u_24u.v(901[10:33])
    wire mco_118;   // mult_24u_24u.v(900[10:17])
    wire mult_24u_24u_0_pp_10_39;   // mult_24u_24u.v(899[10:33])
    wire mult_24u_24u_0_pp_10_40;   // mult_24u_24u.v(898[10:33])
    wire mco_117;   // mult_24u_24u.v(897[10:17])
    wire mult_24u_24u_0_pp_10_37;   // mult_24u_24u.v(896[10:33])
    wire mult_24u_24u_0_pp_10_38;   // mult_24u_24u.v(895[10:33])
    wire mco_116;   // mult_24u_24u.v(894[10:17])
    wire mult_24u_24u_0_pp_10_35;   // mult_24u_24u.v(893[10:33])
    wire mult_24u_24u_0_pp_10_36;   // mult_24u_24u.v(892[10:33])
    wire mco_115;   // mult_24u_24u.v(891[10:17])
    wire mult_24u_24u_0_pp_10_33;   // mult_24u_24u.v(890[10:33])
    wire mult_24u_24u_0_pp_10_34;   // mult_24u_24u.v(889[10:33])
    wire mco_114;   // mult_24u_24u.v(888[10:17])
    wire mult_24u_24u_0_pp_10_31;   // mult_24u_24u.v(887[10:33])
    wire mult_24u_24u_0_pp_10_32;   // mult_24u_24u.v(886[10:33])
    wire mco_113;   // mult_24u_24u.v(885[10:17])
    wire mult_24u_24u_0_pp_10_29;   // mult_24u_24u.v(884[10:33])
    wire mult_24u_24u_0_pp_10_30;   // mult_24u_24u.v(883[10:33])
    wire mco_112;   // mult_24u_24u.v(882[10:17])
    wire mult_24u_24u_0_pp_10_27;   // mult_24u_24u.v(881[10:33])
    wire mult_24u_24u_0_pp_10_28;   // mult_24u_24u.v(880[10:33])
    wire mco_111;   // mult_24u_24u.v(879[10:17])
    wire mult_24u_24u_0_pp_10_25;   // mult_24u_24u.v(878[10:33])
    wire mult_24u_24u_0_pp_10_26;   // mult_24u_24u.v(877[10:33])
    wire mco_110;   // mult_24u_24u.v(876[10:17])
    wire mult_24u_24u_0_pp_10_23;   // mult_24u_24u.v(875[10:33])
    wire mult_24u_24u_0_pp_10_24;   // mult_24u_24u.v(874[10:33])
    wire mult_24u_24u_0_cin_lr_20;   // mult_24u_24u.v(873[10:34])
    wire mult_24u_24u_0_pp_10_21;   // mult_24u_24u.v(872[10:33])
    wire mult_24u_24u_0_pp_10_22;   // mult_24u_24u.v(871[10:33])
    wire mco_109;   // mult_24u_24u.v(870[10:17])
    wire mult_24u_24u_0_pp_9_41;   // mult_24u_24u.v(869[10:32])
    wire mult_24u_24u_0_pp_9_42;   // mult_24u_24u.v(868[10:32])
    wire mfco_9;   // mult_24u_24u.v(867[10:16])
    wire mco_108;   // mult_24u_24u.v(866[10:17])
    wire mult_24u_24u_0_pp_9_39;   // mult_24u_24u.v(865[10:32])
    wire mult_24u_24u_0_pp_9_40;   // mult_24u_24u.v(864[10:32])
    wire mco_107;   // mult_24u_24u.v(863[10:17])
    wire mult_24u_24u_0_pp_9_37;   // mult_24u_24u.v(862[10:32])
    wire mult_24u_24u_0_pp_9_38;   // mult_24u_24u.v(861[10:32])
    wire mco_106;   // mult_24u_24u.v(860[10:17])
    wire mult_24u_24u_0_pp_9_35;   // mult_24u_24u.v(859[10:32])
    wire mult_24u_24u_0_pp_9_36;   // mult_24u_24u.v(858[10:32])
    wire mco_105;   // mult_24u_24u.v(857[10:17])
    wire mult_24u_24u_0_pp_9_33;   // mult_24u_24u.v(856[10:32])
    wire mult_24u_24u_0_pp_9_34;   // mult_24u_24u.v(855[10:32])
    wire mco_104;   // mult_24u_24u.v(854[10:17])
    wire mult_24u_24u_0_pp_9_31;   // mult_24u_24u.v(853[10:32])
    wire mult_24u_24u_0_pp_9_32;   // mult_24u_24u.v(852[10:32])
    wire mco_103;   // mult_24u_24u.v(851[10:17])
    wire mult_24u_24u_0_pp_9_29;   // mult_24u_24u.v(850[10:32])
    wire mult_24u_24u_0_pp_9_30;   // mult_24u_24u.v(849[10:32])
    wire mco_102;   // mult_24u_24u.v(848[10:17])
    wire mult_24u_24u_0_pp_9_27;   // mult_24u_24u.v(847[10:32])
    wire mult_24u_24u_0_pp_9_28;   // mult_24u_24u.v(846[10:32])
    wire mco_101;   // mult_24u_24u.v(845[10:17])
    wire mult_24u_24u_0_pp_9_25;   // mult_24u_24u.v(844[10:32])
    wire mult_24u_24u_0_pp_9_26;   // mult_24u_24u.v(843[10:32])
    wire mco_100;   // mult_24u_24u.v(842[10:17])
    wire mult_24u_24u_0_pp_9_23;   // mult_24u_24u.v(841[10:32])
    wire mult_24u_24u_0_pp_9_24;   // mult_24u_24u.v(840[10:32])
    wire mco_99;   // mult_24u_24u.v(839[10:16])
    wire mult_24u_24u_0_pp_9_21;   // mult_24u_24u.v(838[10:32])
    wire mult_24u_24u_0_pp_9_22;   // mult_24u_24u.v(837[10:32])
    wire mult_24u_24u_0_cin_lr_18;   // mult_24u_24u.v(836[10:34])
    wire mult_24u_24u_0_pp_9_19;   // mult_24u_24u.v(835[10:32])
    wire mult_24u_24u_0_pp_9_20;   // mult_24u_24u.v(834[10:32])
    wire mco_98;   // mult_24u_24u.v(833[10:16])
    wire mult_24u_24u_0_pp_8_39;   // mult_24u_24u.v(832[10:32])
    wire mult_24u_24u_0_pp_8_40;   // mult_24u_24u.v(831[10:32])
    wire mfco_8;   // mult_24u_24u.v(830[10:16])
    wire mco_97;   // mult_24u_24u.v(829[10:16])
    wire mult_24u_24u_0_pp_8_37;   // mult_24u_24u.v(828[10:32])
    wire mult_24u_24u_0_pp_8_38;   // mult_24u_24u.v(827[10:32])
    wire mco_96;   // mult_24u_24u.v(826[10:16])
    wire mult_24u_24u_0_pp_8_35;   // mult_24u_24u.v(825[10:32])
    wire mult_24u_24u_0_pp_8_36;   // mult_24u_24u.v(824[10:32])
    wire mco_95;   // mult_24u_24u.v(823[10:16])
    wire mult_24u_24u_0_pp_8_33;   // mult_24u_24u.v(822[10:32])
    wire mult_24u_24u_0_pp_8_34;   // mult_24u_24u.v(821[10:32])
    wire [4:0]n2889;   // mult_3u_2u.v(11[23:24])
    wire [4:0]n3044;   // mult_2u_3u.v(11[23:24])
    wire mco_94;   // mult_24u_24u.v(820[10:16])
    wire mult_24u_24u_0_pp_8_31;   // mult_24u_24u.v(819[10:32])
    wire mult_24u_24u_0_pp_8_32;   // mult_24u_24u.v(818[10:32])
    wire mco_93;   // mult_24u_24u.v(817[10:16])
    wire mult_24u_24u_0_pp_8_29;   // mult_24u_24u.v(816[10:32])
    wire mult_24u_24u_0_pp_8_30;   // mult_24u_24u.v(815[10:32])
    wire mco_92;   // mult_24u_24u.v(814[10:16])
    wire mult_24u_24u_0_pp_8_27;   // mult_24u_24u.v(813[10:32])
    wire mult_24u_24u_0_pp_8_28;   // mult_24u_24u.v(812[10:32])
    wire mco_91;   // mult_24u_24u.v(811[10:16])
    wire mult_24u_24u_0_pp_8_25;   // mult_24u_24u.v(810[10:32])
    wire mult_24u_24u_0_pp_8_26;   // mult_24u_24u.v(809[10:32])
    wire mco_90;   // mult_24u_24u.v(808[10:16])
    wire mult_24u_24u_0_pp_8_23;   // mult_24u_24u.v(807[10:32])
    wire mult_24u_24u_0_pp_8_24;   // mult_24u_24u.v(806[10:32])
    wire mco_89;   // mult_24u_24u.v(805[10:16])
    wire mult_24u_24u_0_pp_8_21;   // mult_24u_24u.v(804[10:32])
    wire mult_24u_24u_0_pp_8_22;   // mult_24u_24u.v(803[10:32])
    wire mco_88;   // mult_24u_24u.v(802[10:16])
    wire mult_24u_24u_0_pp_8_19;   // mult_24u_24u.v(801[10:32])
    wire mult_24u_24u_0_pp_8_20;   // mult_24u_24u.v(800[10:32])
    wire mult_24u_24u_0_cin_lr_16;   // mult_24u_24u.v(799[10:34])
    wire mult_24u_24u_0_pp_8_17;   // mult_24u_24u.v(798[10:32])
    wire mult_24u_24u_0_pp_8_18;   // mult_24u_24u.v(797[10:32])
    wire mco_87;   // mult_24u_24u.v(796[10:16])
    wire mult_24u_24u_0_pp_7_37;   // mult_24u_24u.v(795[10:32])
    wire mult_24u_24u_0_pp_7_38;   // mult_24u_24u.v(794[10:32])
    wire mfco_7;   // mult_24u_24u.v(793[10:16])
    wire mco_86;   // mult_24u_24u.v(792[10:16])
    wire mult_24u_24u_0_pp_7_35;   // mult_24u_24u.v(791[10:32])
    wire mult_24u_24u_0_pp_7_36;   // mult_24u_24u.v(790[10:32])
    wire mco_85;   // mult_24u_24u.v(789[10:16])
    wire mult_24u_24u_0_pp_7_33;   // mult_24u_24u.v(788[10:32])
    wire mult_24u_24u_0_pp_7_34;   // mult_24u_24u.v(787[10:32])
    wire mco_84;   // mult_24u_24u.v(786[10:16])
    wire mult_24u_24u_0_pp_7_31;   // mult_24u_24u.v(785[10:32])
    wire mult_24u_24u_0_pp_7_32;   // mult_24u_24u.v(784[10:32])
    wire mco_83;   // mult_24u_24u.v(783[10:16])
    wire mult_24u_24u_0_pp_7_29;   // mult_24u_24u.v(782[10:32])
    wire mult_24u_24u_0_pp_7_30;   // mult_24u_24u.v(781[10:32])
    wire mco_82;   // mult_24u_24u.v(780[10:16])
    wire mult_24u_24u_0_pp_7_27;   // mult_24u_24u.v(779[10:32])
    wire mult_24u_24u_0_pp_7_28;   // mult_24u_24u.v(778[10:32])
    wire mco_81;   // mult_24u_24u.v(777[10:16])
    wire mult_24u_24u_0_pp_7_25;   // mult_24u_24u.v(776[10:32])
    wire mult_24u_24u_0_pp_7_26;   // mult_24u_24u.v(775[10:32])
    wire mco_80;   // mult_24u_24u.v(774[10:16])
    wire mult_24u_24u_0_pp_7_23;   // mult_24u_24u.v(773[10:32])
    wire mult_24u_24u_0_pp_7_24;   // mult_24u_24u.v(772[10:32])
    wire mco_79;   // mult_24u_24u.v(771[10:16])
    wire mult_24u_24u_0_pp_7_21;   // mult_24u_24u.v(770[10:32])
    wire mult_24u_24u_0_pp_7_22;   // mult_24u_24u.v(769[10:32])
    wire mco_78;   // mult_24u_24u.v(768[10:16])
    wire mult_24u_24u_0_pp_7_19;   // mult_24u_24u.v(767[10:32])
    wire mult_24u_24u_0_pp_7_20;   // mult_24u_24u.v(766[10:32])
    wire mco_77;   // mult_24u_24u.v(765[10:16])
    wire mult_24u_24u_0_pp_7_17;   // mult_24u_24u.v(764[10:32])
    wire mult_24u_24u_0_pp_7_18;   // mult_24u_24u.v(763[10:32])
    wire mult_24u_24u_0_cin_lr_14;   // mult_24u_24u.v(762[10:34])
    wire mult_24u_24u_0_pp_7_15;   // mult_24u_24u.v(761[10:32])
    wire mult_24u_24u_0_pp_7_16;   // mult_24u_24u.v(760[10:32])
    wire mco_76;   // mult_24u_24u.v(759[10:16])
    wire mult_24u_24u_0_pp_6_35;   // mult_24u_24u.v(758[10:32])
    wire mult_24u_24u_0_pp_6_36;   // mult_24u_24u.v(757[10:32])
    wire mfco_6;   // mult_24u_24u.v(756[10:16])
    wire mco_75;   // mult_24u_24u.v(755[10:16])
    wire mult_24u_24u_0_pp_6_33;   // mult_24u_24u.v(754[10:32])
    wire mult_24u_24u_0_pp_6_34;   // mult_24u_24u.v(753[10:32])
    wire mco_74;   // mult_24u_24u.v(752[10:16])
    wire mult_24u_24u_0_pp_6_31;   // mult_24u_24u.v(751[10:32])
    wire mult_24u_24u_0_pp_6_32;   // mult_24u_24u.v(750[10:32])
    wire mco_73;   // mult_24u_24u.v(749[10:16])
    wire mult_24u_24u_0_pp_6_29;   // mult_24u_24u.v(748[10:32])
    wire mult_24u_24u_0_pp_6_30;   // mult_24u_24u.v(747[10:32])
    wire mco_72;   // mult_24u_24u.v(746[10:16])
    wire mult_24u_24u_0_pp_6_27;   // mult_24u_24u.v(745[10:32])
    wire mult_24u_24u_0_pp_6_28;   // mult_24u_24u.v(744[10:32])
    wire mco_71;   // mult_24u_24u.v(743[10:16])
    wire mult_24u_24u_0_pp_6_25;   // mult_24u_24u.v(742[10:32])
    wire mult_24u_24u_0_pp_6_26;   // mult_24u_24u.v(741[10:32])
    wire mco_70;   // mult_24u_24u.v(740[10:16])
    wire mult_24u_24u_0_pp_6_23;   // mult_24u_24u.v(739[10:32])
    wire mult_24u_24u_0_pp_6_24;   // mult_24u_24u.v(738[10:32])
    wire mco_69;   // mult_24u_24u.v(737[10:16])
    wire mult_24u_24u_0_pp_6_21;   // mult_24u_24u.v(736[10:32])
    wire mult_24u_24u_0_pp_6_22;   // mult_24u_24u.v(735[10:32])
    wire mco_68;   // mult_24u_24u.v(734[10:16])
    wire mult_24u_24u_0_pp_6_19;   // mult_24u_24u.v(733[10:32])
    wire mult_24u_24u_0_pp_6_20;   // mult_24u_24u.v(732[10:32])
    wire mco_67;   // mult_24u_24u.v(731[10:16])
    wire mult_24u_24u_0_pp_6_17;   // mult_24u_24u.v(730[10:32])
    wire mult_24u_24u_0_pp_6_18;   // mult_24u_24u.v(729[10:32])
    wire mco_66;   // mult_24u_24u.v(728[10:16])
    wire mult_24u_24u_0_pp_6_15;   // mult_24u_24u.v(727[10:32])
    wire mult_24u_24u_0_pp_6_16;   // mult_24u_24u.v(726[10:32])
    wire mult_24u_24u_0_cin_lr_12;   // mult_24u_24u.v(725[10:34])
    wire mult_24u_24u_0_pp_6_13;   // mult_24u_24u.v(724[10:32])
    wire mult_24u_24u_0_pp_6_14;   // mult_24u_24u.v(723[10:32])
    wire mco_65;   // mult_24u_24u.v(722[10:16])
    wire mult_24u_24u_0_pp_5_33;   // mult_24u_24u.v(721[10:32])
    wire mult_24u_24u_0_pp_5_34;   // mult_24u_24u.v(720[10:32])
    wire mfco_5;   // mult_24u_24u.v(719[10:16])
    wire mco_64;   // mult_24u_24u.v(718[10:16])
    wire mult_24u_24u_0_pp_5_31;   // mult_24u_24u.v(717[10:32])
    wire mult_24u_24u_0_pp_5_32;   // mult_24u_24u.v(716[10:32])
    wire mco_63;   // mult_24u_24u.v(715[10:16])
    wire mult_24u_24u_0_pp_5_29;   // mult_24u_24u.v(714[10:32])
    wire mult_24u_24u_0_pp_5_30;   // mult_24u_24u.v(713[10:32])
    wire mco_62;   // mult_24u_24u.v(712[10:16])
    wire mult_24u_24u_0_pp_5_27;   // mult_24u_24u.v(711[10:32])
    wire mult_24u_24u_0_pp_5_28;   // mult_24u_24u.v(710[10:32])
    wire mco_61;   // mult_24u_24u.v(709[10:16])
    wire mult_24u_24u_0_pp_5_25;   // mult_24u_24u.v(708[10:32])
    wire mult_24u_24u_0_pp_5_26;   // mult_24u_24u.v(707[10:32])
    wire mco_60;   // mult_24u_24u.v(706[10:16])
    wire mult_24u_24u_0_pp_5_23;   // mult_24u_24u.v(705[10:32])
    wire mult_24u_24u_0_pp_5_24;   // mult_24u_24u.v(704[10:32])
    wire mco_59;   // mult_24u_24u.v(703[10:16])
    wire mult_24u_24u_0_pp_5_21;   // mult_24u_24u.v(702[10:32])
    wire mult_24u_24u_0_pp_5_22;   // mult_24u_24u.v(701[10:32])
    wire mco_58;   // mult_24u_24u.v(700[10:16])
    wire mult_24u_24u_0_pp_5_19;   // mult_24u_24u.v(699[10:32])
    wire mult_24u_24u_0_pp_5_20;   // mult_24u_24u.v(698[10:32])
    wire mco_57;   // mult_24u_24u.v(697[10:16])
    wire mult_24u_24u_0_pp_5_17;   // mult_24u_24u.v(696[10:32])
    wire mult_24u_24u_0_pp_5_18;   // mult_24u_24u.v(695[10:32])
    wire mco_56;   // mult_24u_24u.v(694[10:16])
    wire mult_24u_24u_0_pp_5_15;   // mult_24u_24u.v(693[10:32])
    wire mult_24u_24u_0_pp_5_16;   // mult_24u_24u.v(692[10:32])
    wire mco_55;   // mult_24u_24u.v(691[10:16])
    wire mult_24u_24u_0_pp_5_13;   // mult_24u_24u.v(690[10:32])
    wire mult_24u_24u_0_pp_5_14;   // mult_24u_24u.v(689[10:32])
    wire mult_24u_24u_0_cin_lr_10;   // mult_24u_24u.v(688[10:34])
    wire mult_24u_24u_0_pp_5_11;   // mult_24u_24u.v(687[10:32])
    wire mult_24u_24u_0_pp_5_12;   // mult_24u_24u.v(686[10:32])
    wire mco_54;   // mult_24u_24u.v(685[10:16])
    wire mult_24u_24u_0_pp_4_31;   // mult_24u_24u.v(684[10:32])
    wire mult_24u_24u_0_pp_4_32;   // mult_24u_24u.v(683[10:32])
    wire mfco_4;   // mult_24u_24u.v(682[10:16])
    wire mco_53;   // mult_24u_24u.v(681[10:16])
    wire mult_24u_24u_0_pp_4_29;   // mult_24u_24u.v(680[10:32])
    wire mult_24u_24u_0_pp_4_30;   // mult_24u_24u.v(679[10:32])
    wire mco_52;   // mult_24u_24u.v(678[10:16])
    wire mult_24u_24u_0_pp_4_27;   // mult_24u_24u.v(677[10:32])
    wire mult_24u_24u_0_pp_4_28;   // mult_24u_24u.v(676[10:32])
    wire mco_51;   // mult_24u_24u.v(675[10:16])
    wire mult_24u_24u_0_pp_4_25;   // mult_24u_24u.v(674[10:32])
    wire mult_24u_24u_0_pp_4_26;   // mult_24u_24u.v(673[10:32])
    wire mco_50;   // mult_24u_24u.v(672[10:16])
    wire mult_24u_24u_0_pp_4_23;   // mult_24u_24u.v(671[10:32])
    wire mult_24u_24u_0_pp_4_24;   // mult_24u_24u.v(670[10:32])
    wire mco_49;   // mult_24u_24u.v(669[10:16])
    wire mult_24u_24u_0_pp_4_21;   // mult_24u_24u.v(668[10:32])
    wire mult_24u_24u_0_pp_4_22;   // mult_24u_24u.v(667[10:32])
    wire mco_48;   // mult_24u_24u.v(666[10:16])
    wire mult_24u_24u_0_pp_4_19;   // mult_24u_24u.v(665[10:32])
    wire mult_24u_24u_0_pp_4_20;   // mult_24u_24u.v(664[10:32])
    wire mco_47;   // mult_24u_24u.v(663[10:16])
    wire mult_24u_24u_0_pp_4_17;   // mult_24u_24u.v(662[10:32])
    wire mult_24u_24u_0_pp_4_18;   // mult_24u_24u.v(661[10:32])
    wire mco_46;   // mult_24u_24u.v(660[10:16])
    wire mult_24u_24u_0_pp_4_15;   // mult_24u_24u.v(659[10:32])
    wire mult_24u_24u_0_pp_4_16;   // mult_24u_24u.v(658[10:32])
    wire mco_45;   // mult_24u_24u.v(657[10:16])
    wire mult_24u_24u_0_pp_4_13;   // mult_24u_24u.v(656[10:32])
    wire mult_24u_24u_0_pp_4_14;   // mult_24u_24u.v(655[10:32])
    wire mco_44;   // mult_24u_24u.v(654[10:16])
    wire mult_24u_24u_0_pp_4_11;   // mult_24u_24u.v(653[10:32])
    wire mult_24u_24u_0_pp_4_12;   // mult_24u_24u.v(652[10:32])
    wire mult_24u_24u_0_cin_lr_8;   // mult_24u_24u.v(651[10:33])
    wire mult_24u_24u_0_pp_4_9;   // mult_24u_24u.v(650[10:31])
    wire mult_24u_24u_0_pp_4_10;   // mult_24u_24u.v(649[10:32])
    wire mco_43;   // mult_24u_24u.v(648[10:16])
    wire mult_24u_24u_0_pp_3_29;   // mult_24u_24u.v(647[10:32])
    wire mult_24u_24u_0_pp_3_30;   // mult_24u_24u.v(646[10:32])
    wire mfco_3;   // mult_24u_24u.v(645[10:16])
    wire mco_42;   // mult_24u_24u.v(644[10:16])
    wire mult_24u_24u_0_pp_3_27;   // mult_24u_24u.v(643[10:32])
    wire mult_24u_24u_0_pp_3_28;   // mult_24u_24u.v(642[10:32])
    wire mco_41;   // mult_24u_24u.v(641[10:16])
    wire mult_24u_24u_0_pp_3_25;   // mult_24u_24u.v(640[10:32])
    wire mult_24u_24u_0_pp_3_26;   // mult_24u_24u.v(639[10:32])
    wire mco_40;   // mult_24u_24u.v(638[10:16])
    wire mult_24u_24u_0_pp_3_23;   // mult_24u_24u.v(637[10:32])
    wire mult_24u_24u_0_pp_3_24;   // mult_24u_24u.v(636[10:32])
    wire mco_39;   // mult_24u_24u.v(635[10:16])
    wire mult_24u_24u_0_pp_3_21;   // mult_24u_24u.v(634[10:32])
    wire mult_24u_24u_0_pp_3_22;   // mult_24u_24u.v(633[10:32])
    wire mco_38;   // mult_24u_24u.v(632[10:16])
    wire mult_24u_24u_0_pp_3_19;   // mult_24u_24u.v(631[10:32])
    wire mult_24u_24u_0_pp_3_20;   // mult_24u_24u.v(630[10:32])
    wire mco_37;   // mult_24u_24u.v(629[10:16])
    wire mult_24u_24u_0_pp_3_17;   // mult_24u_24u.v(628[10:32])
    wire mult_24u_24u_0_pp_3_18;   // mult_24u_24u.v(627[10:32])
    wire mco_36;   // mult_24u_24u.v(626[10:16])
    wire mult_24u_24u_0_pp_3_15;   // mult_24u_24u.v(625[10:32])
    wire mult_24u_24u_0_pp_3_16;   // mult_24u_24u.v(624[10:32])
    wire mco_35;   // mult_24u_24u.v(623[10:16])
    wire mult_24u_24u_0_pp_3_13;   // mult_24u_24u.v(622[10:32])
    wire mult_24u_24u_0_pp_3_14;   // mult_24u_24u.v(621[10:32])
    wire mco_34;   // mult_24u_24u.v(620[10:16])
    wire mult_24u_24u_0_pp_3_11;   // mult_24u_24u.v(619[10:32])
    wire mult_24u_24u_0_pp_3_12;   // mult_24u_24u.v(618[10:32])
    wire mco_33;   // mult_24u_24u.v(617[10:16])
    wire mult_24u_24u_0_pp_3_9;   // mult_24u_24u.v(616[10:31])
    wire mult_24u_24u_0_pp_3_10;   // mult_24u_24u.v(615[10:32])
    wire mult_24u_24u_0_cin_lr_6;   // mult_24u_24u.v(614[10:33])
    wire mult_24u_24u_0_pp_3_7;   // mult_24u_24u.v(613[10:31])
    wire mult_24u_24u_0_pp_3_8;   // mult_24u_24u.v(612[10:31])
    wire mco_32;   // mult_24u_24u.v(611[10:16])
    wire mult_24u_24u_0_pp_2_27;   // mult_24u_24u.v(610[10:32])
    wire mult_24u_24u_0_pp_2_28;   // mult_24u_24u.v(609[10:32])
    wire mfco_2;   // mult_24u_24u.v(608[10:16])
    wire mco_31;   // mult_24u_24u.v(607[10:16])
    wire mult_24u_24u_0_pp_2_25;   // mult_24u_24u.v(606[10:32])
    wire mult_24u_24u_0_pp_2_26;   // mult_24u_24u.v(605[10:32])
    wire mco_30;   // mult_24u_24u.v(604[10:16])
    wire mult_24u_24u_0_pp_2_23;   // mult_24u_24u.v(603[10:32])
    wire mult_24u_24u_0_pp_2_24;   // mult_24u_24u.v(602[10:32])
    wire mco_29;   // mult_24u_24u.v(601[10:16])
    wire mult_24u_24u_0_pp_2_21;   // mult_24u_24u.v(600[10:32])
    wire mult_24u_24u_0_pp_2_22;   // mult_24u_24u.v(599[10:32])
    wire mco_28;   // mult_24u_24u.v(598[10:16])
    wire mult_24u_24u_0_pp_2_19;   // mult_24u_24u.v(597[10:32])
    wire mult_24u_24u_0_pp_2_20;   // mult_24u_24u.v(596[10:32])
    wire mco_27;   // mult_24u_24u.v(595[10:16])
    wire mult_24u_24u_0_pp_2_17;   // mult_24u_24u.v(594[10:32])
    wire mult_24u_24u_0_pp_2_18;   // mult_24u_24u.v(593[10:32])
    wire mco_26;   // mult_24u_24u.v(592[10:16])
    wire mult_24u_24u_0_pp_2_15;   // mult_24u_24u.v(591[10:32])
    wire mult_24u_24u_0_pp_2_16;   // mult_24u_24u.v(590[10:32])
    wire mco_25;   // mult_24u_24u.v(589[10:16])
    wire mult_24u_24u_0_pp_2_13;   // mult_24u_24u.v(588[10:32])
    wire mult_24u_24u_0_pp_2_14;   // mult_24u_24u.v(587[10:32])
    wire mco_24;   // mult_24u_24u.v(586[10:16])
    wire mult_24u_24u_0_pp_2_11;   // mult_24u_24u.v(585[10:32])
    wire mult_24u_24u_0_pp_2_12;   // mult_24u_24u.v(584[10:32])
    wire mco_23;   // mult_24u_24u.v(583[10:16])
    wire mult_24u_24u_0_pp_2_9;   // mult_24u_24u.v(582[10:31])
    wire mult_24u_24u_0_pp_2_10;   // mult_24u_24u.v(581[10:32])
    wire mco_22;   // mult_24u_24u.v(580[10:16])
    wire mult_24u_24u_0_pp_2_7;   // mult_24u_24u.v(579[10:31])
    wire mult_24u_24u_0_pp_2_8;   // mult_24u_24u.v(578[10:31])
    wire mult_24u_24u_0_cin_lr_4;   // mult_24u_24u.v(577[10:33])
    wire mult_24u_24u_0_pp_2_5;   // mult_24u_24u.v(576[10:31])
    wire mult_24u_24u_0_pp_2_6;   // mult_24u_24u.v(575[10:31])
    wire mco_21;   // mult_24u_24u.v(574[10:16])
    wire mult_24u_24u_0_pp_1_25;   // mult_24u_24u.v(573[10:32])
    wire mult_24u_24u_0_pp_1_26;   // mult_24u_24u.v(572[10:32])
    wire mfco_1;   // mult_24u_24u.v(571[10:16])
    wire mco_20;   // mult_24u_24u.v(570[10:16])
    wire mult_24u_24u_0_pp_1_23;   // mult_24u_24u.v(569[10:32])
    wire mult_24u_24u_0_pp_1_24;   // mult_24u_24u.v(568[10:32])
    wire mco_19;   // mult_24u_24u.v(567[10:16])
    wire mult_24u_24u_0_pp_1_21;   // mult_24u_24u.v(566[10:32])
    wire mult_24u_24u_0_pp_1_22;   // mult_24u_24u.v(565[10:32])
    wire mco_18;   // mult_24u_24u.v(564[10:16])
    wire mult_24u_24u_0_pp_1_19;   // mult_24u_24u.v(563[10:32])
    wire mult_24u_24u_0_pp_1_20;   // mult_24u_24u.v(562[10:32])
    wire mco_17;   // mult_24u_24u.v(561[10:16])
    wire mult_24u_24u_0_pp_1_17;   // mult_24u_24u.v(560[10:32])
    wire mult_24u_24u_0_pp_1_18;   // mult_24u_24u.v(559[10:32])
    wire mco_16;   // mult_24u_24u.v(558[10:16])
    wire mult_24u_24u_0_pp_1_15;   // mult_24u_24u.v(557[10:32])
    wire mult_24u_24u_0_pp_1_16;   // mult_24u_24u.v(556[10:32])
    wire mco_15;   // mult_24u_24u.v(555[10:16])
    wire mult_24u_24u_0_pp_1_13;   // mult_24u_24u.v(554[10:32])
    wire mult_24u_24u_0_pp_1_14;   // mult_24u_24u.v(553[10:32])
    wire mco_14;   // mult_24u_24u.v(552[10:16])
    wire mult_24u_24u_0_pp_1_11;   // mult_24u_24u.v(551[10:32])
    wire mult_24u_24u_0_pp_1_12;   // mult_24u_24u.v(550[10:32])
    wire mco_13;   // mult_24u_24u.v(549[10:16])
    wire mult_24u_24u_0_pp_1_9;   // mult_24u_24u.v(548[10:31])
    wire mult_24u_24u_0_pp_1_10;   // mult_24u_24u.v(547[10:32])
    wire mco_12;   // mult_24u_24u.v(546[10:16])
    wire mult_24u_24u_0_pp_1_7;   // mult_24u_24u.v(545[10:31])
    wire mult_24u_24u_0_pp_1_8;   // mult_24u_24u.v(544[10:31])
    wire mco_11;   // mult_24u_24u.v(543[10:16])
    wire mult_24u_24u_0_pp_1_5;   // mult_24u_24u.v(542[10:31])
    wire mult_24u_24u_0_pp_1_6;   // mult_24u_24u.v(541[10:31])
    wire mult_24u_24u_0_cin_lr_2;   // mult_24u_24u.v(540[10:33])
    wire mult_24u_24u_0_pp_1_3;   // mult_24u_24u.v(539[10:31])
    wire mult_24u_24u_0_pp_1_4;   // mult_24u_24u.v(538[10:31])
    wire mco_10;   // mult_24u_24u.v(537[10:16])
    wire mult_24u_24u_0_pp_0_23;   // mult_24u_24u.v(536[10:32])
    wire mult_24u_24u_0_pp_0_24;   // mult_24u_24u.v(535[10:32])
    wire mfco;   // mult_24u_24u.v(534[10:14])
    wire mco_9;   // mult_24u_24u.v(533[10:15])
    wire mult_24u_24u_0_pp_0_21;   // mult_24u_24u.v(532[10:32])
    wire mult_24u_24u_0_pp_0_22;   // mult_24u_24u.v(531[10:32])
    wire mco_8;   // mult_24u_24u.v(530[10:15])
    wire mult_24u_24u_0_pp_0_19;   // mult_24u_24u.v(529[10:32])
    wire mult_24u_24u_0_pp_0_20;   // mult_24u_24u.v(528[10:32])
    wire mco_7;   // mult_24u_24u.v(527[10:15])
    wire mult_24u_24u_0_pp_0_17;   // mult_24u_24u.v(526[10:32])
    wire mult_24u_24u_0_pp_0_18;   // mult_24u_24u.v(525[10:32])
    wire mco_6;   // mult_24u_24u.v(524[10:15])
    wire mult_24u_24u_0_pp_0_15;   // mult_24u_24u.v(523[10:32])
    wire mult_24u_24u_0_pp_0_16;   // mult_24u_24u.v(522[10:32])
    wire mco_5;   // mult_24u_24u.v(521[10:15])
    wire mult_24u_24u_0_pp_0_13;   // mult_24u_24u.v(520[10:32])
    wire mult_24u_24u_0_pp_0_14;   // mult_24u_24u.v(519[10:32])
    wire mco_4;   // mult_24u_24u.v(518[10:15])
    wire mult_24u_24u_0_pp_0_11;   // mult_24u_24u.v(517[10:32])
    wire mult_24u_24u_0_pp_0_12;   // mult_24u_24u.v(516[10:32])
    wire mco_3;   // mult_24u_24u.v(515[10:15])
    wire mult_24u_24u_0_pp_0_9;   // mult_24u_24u.v(514[10:31])
    wire mult_24u_24u_0_pp_0_10;   // mult_24u_24u.v(513[10:32])
    wire mco_2;   // mult_24u_24u.v(512[10:15])
    wire mult_24u_24u_0_pp_0_7;   // mult_24u_24u.v(511[10:31])
    wire mult_24u_24u_0_pp_0_8;   // mult_24u_24u.v(510[10:31])
    wire mco_1;   // mult_24u_24u.v(509[10:15])
    wire mult_24u_24u_0_pp_0_5;   // mult_24u_24u.v(508[10:31])
    wire mult_24u_24u_0_pp_0_6;   // mult_24u_24u.v(507[10:31])
    wire mco;   // mult_24u_24u.v(506[10:13])
    wire mult_24u_24u_0_pp_0_3;   // mult_24u_24u.v(505[10:31])
    wire mult_24u_24u_0_pp_0_4;   // mult_24u_24u.v(504[10:31])
    wire mult_24u_24u_0_cin_lr_0;   // mult_24u_24u.v(503[10:33])
    wire mult_24u_24u_0_pp_0_2;   // mult_24u_24u.v(501[10:31])
    wire s_mult_24u_24u_0_8_47;   // mult_24u_24u.v(500[10:31])
    wire co_t_mult_24u_24u_0_10_16;   // mult_24u_24u.v(499[10:35])
    wire s_mult_24u_24u_0_9_45;   // mult_24u_24u.v(497[10:31])
    wire s_mult_24u_24u_0_8_46;   // mult_24u_24u.v(496[10:31])
    wire s_mult_24u_24u_0_8_45;   // mult_24u_24u.v(495[10:31])
    wire co_t_mult_24u_24u_0_10_15;   // mult_24u_24u.v(494[10:35])
    wire s_mult_24u_24u_0_9_44;   // mult_24u_24u.v(493[10:31])
    wire s_mult_24u_24u_0_9_43;   // mult_24u_24u.v(492[10:31])
    wire s_mult_24u_24u_0_8_44;   // mult_24u_24u.v(491[10:31])
    wire s_mult_24u_24u_0_8_43;   // mult_24u_24u.v(490[10:31])
    wire co_t_mult_24u_24u_0_10_14;   // mult_24u_24u.v(489[10:35])
    wire s_mult_24u_24u_0_9_42;   // mult_24u_24u.v(488[10:31])
    wire s_mult_24u_24u_0_9_41;   // mult_24u_24u.v(487[10:31])
    wire s_mult_24u_24u_0_8_42;   // mult_24u_24u.v(486[10:31])
    wire s_mult_24u_24u_0_8_41;   // mult_24u_24u.v(485[10:31])
    wire co_t_mult_24u_24u_0_10_13;   // mult_24u_24u.v(484[10:35])
    wire s_mult_24u_24u_0_9_40;   // mult_24u_24u.v(483[10:31])
    wire s_mult_24u_24u_0_9_39;   // mult_24u_24u.v(482[10:31])
    wire s_mult_24u_24u_0_8_40;   // mult_24u_24u.v(481[10:31])
    wire s_mult_24u_24u_0_8_39;   // mult_24u_24u.v(480[10:31])
    wire co_t_mult_24u_24u_0_10_12;   // mult_24u_24u.v(479[10:35])
    wire s_mult_24u_24u_0_9_38;   // mult_24u_24u.v(478[10:31])
    wire s_mult_24u_24u_0_9_37;   // mult_24u_24u.v(477[10:31])
    wire s_mult_24u_24u_0_8_38;   // mult_24u_24u.v(476[10:31])
    wire s_mult_24u_24u_0_8_37;   // mult_24u_24u.v(475[10:31])
    wire co_t_mult_24u_24u_0_10_11;   // mult_24u_24u.v(474[10:35])
    wire s_mult_24u_24u_0_9_36;   // mult_24u_24u.v(473[10:31])
    wire s_mult_24u_24u_0_9_35;   // mult_24u_24u.v(472[10:31])
    wire s_mult_24u_24u_0_8_36;   // mult_24u_24u.v(471[10:31])
    wire s_mult_24u_24u_0_8_35;   // mult_24u_24u.v(470[10:31])
    wire co_t_mult_24u_24u_0_10_10;   // mult_24u_24u.v(469[10:35])
    wire s_mult_24u_24u_0_9_34;   // mult_24u_24u.v(468[10:31])
    wire s_mult_24u_24u_0_9_33;   // mult_24u_24u.v(467[10:31])
    wire s_mult_24u_24u_0_8_34;   // mult_24u_24u.v(466[10:31])
    wire s_mult_24u_24u_0_8_33;   // mult_24u_24u.v(465[10:31])
    wire co_t_mult_24u_24u_0_10_9;   // mult_24u_24u.v(464[10:34])
    wire s_mult_24u_24u_0_9_32;   // mult_24u_24u.v(463[10:31])
    wire s_mult_24u_24u_0_9_31;   // mult_24u_24u.v(462[10:31])
    wire s_mult_24u_24u_0_8_32;   // mult_24u_24u.v(461[10:31])
    wire s_mult_24u_24u_0_8_31;   // mult_24u_24u.v(460[10:31])
    wire co_t_mult_24u_24u_0_10_8;   // mult_24u_24u.v(459[10:34])
    wire s_mult_24u_24u_0_9_30;   // mult_24u_24u.v(458[10:31])
    wire s_mult_24u_24u_0_9_29;   // mult_24u_24u.v(457[10:31])
    wire s_mult_24u_24u_0_8_30;   // mult_24u_24u.v(456[10:31])
    wire s_mult_24u_24u_0_8_29;   // mult_24u_24u.v(455[10:31])
    wire co_t_mult_24u_24u_0_10_7;   // mult_24u_24u.v(454[10:34])
    wire s_mult_24u_24u_0_9_28;   // mult_24u_24u.v(453[10:31])
    wire s_mult_24u_24u_0_9_27;   // mult_24u_24u.v(452[10:31])
    wire s_mult_24u_24u_0_8_28;   // mult_24u_24u.v(451[10:31])
    wire s_mult_24u_24u_0_8_27;   // mult_24u_24u.v(450[10:31])
    wire co_t_mult_24u_24u_0_10_6;   // mult_24u_24u.v(449[10:34])
    wire s_mult_24u_24u_0_9_26;   // mult_24u_24u.v(448[10:31])
    wire s_mult_24u_24u_0_9_25;   // mult_24u_24u.v(447[10:31])
    wire s_mult_24u_24u_0_8_26;   // mult_24u_24u.v(446[10:31])
    wire s_mult_24u_24u_0_8_25;   // mult_24u_24u.v(445[10:31])
    wire co_t_mult_24u_24u_0_10_5;   // mult_24u_24u.v(444[10:34])
    wire s_mult_24u_24u_0_9_24;   // mult_24u_24u.v(443[10:31])
    wire s_mult_24u_24u_0_9_23;   // mult_24u_24u.v(442[10:31])
    wire s_mult_24u_24u_0_8_24;   // mult_24u_24u.v(441[10:31])
    wire s_mult_24u_24u_0_8_23;   // mult_24u_24u.v(440[10:31])
    wire co_t_mult_24u_24u_0_10_4;   // mult_24u_24u.v(439[10:34])
    wire s_mult_24u_24u_0_9_22;   // mult_24u_24u.v(438[10:31])
    wire s_mult_24u_24u_0_9_21;   // mult_24u_24u.v(437[10:31])
    wire s_mult_24u_24u_0_8_22;   // mult_24u_24u.v(436[10:31])
    wire s_mult_24u_24u_0_8_21;   // mult_24u_24u.v(435[10:31])
    wire co_t_mult_24u_24u_0_10_3;   // mult_24u_24u.v(434[10:34])
    wire s_mult_24u_24u_0_9_20;   // mult_24u_24u.v(433[10:31])
    wire s_mult_24u_24u_0_9_19;   // mult_24u_24u.v(432[10:31])
    wire s_mult_24u_24u_0_8_20;   // mult_24u_24u.v(431[10:31])
    wire s_mult_24u_24u_0_4_19;   // mult_24u_24u.v(430[10:31])
    wire co_t_mult_24u_24u_0_10_2;   // mult_24u_24u.v(429[10:34])
    wire s_mult_24u_24u_0_9_18;   // mult_24u_24u.v(428[10:31])
    wire s_mult_24u_24u_0_9_17;   // mult_24u_24u.v(427[10:31])
    wire s_mult_24u_24u_0_4_18;   // mult_24u_24u.v(426[10:31])
    wire co_t_mult_24u_24u_0_10_1;   // mult_24u_24u.v(425[10:34])
    wire s_mult_24u_24u_0_9_16;   // mult_24u_24u.v(424[10:31])
    wire mult_24u_24u_0_pp_8_16;   // mult_24u_24u.v(423[10:32])
    wire co_mult_24u_24u_0_9_19;   // mult_24u_24u.v(422[10:32])
    wire s_mult_24u_24u_0_7_43;   // mult_24u_24u.v(421[10:31])
    wire co_mult_24u_24u_0_9_18;   // mult_24u_24u.v(420[10:32])
    wire s_mult_24u_24u_0_7_42;   // mult_24u_24u.v(419[10:31])
    wire s_mult_24u_24u_0_7_41;   // mult_24u_24u.v(418[10:31])
    wire co_mult_24u_24u_0_9_17;   // mult_24u_24u.v(417[10:32])
    wire s_mult_24u_24u_0_7_40;   // mult_24u_24u.v(416[10:31])
    wire s_mult_24u_24u_0_7_39;   // mult_24u_24u.v(415[10:31])
    wire co_mult_24u_24u_0_9_16;   // mult_24u_24u.v(414[10:32])
    wire s_mult_24u_24u_0_7_38;   // mult_24u_24u.v(413[10:31])
    wire s_mult_24u_24u_0_7_37;   // mult_24u_24u.v(412[10:31])
    wire co_mult_24u_24u_0_9_15;   // mult_24u_24u.v(411[10:32])
    wire s_mult_24u_24u_0_6_35;   // mult_24u_24u.v(410[10:31])
    wire s_mult_24u_24u_0_7_36;   // mult_24u_24u.v(409[10:31])
    wire s_mult_24u_24u_0_7_35;   // mult_24u_24u.v(408[10:31])
    wire co_mult_24u_24u_0_9_14;   // mult_24u_24u.v(407[10:32])
    wire s_mult_24u_24u_0_6_34;   // mult_24u_24u.v(406[10:31])
    wire s_mult_24u_24u_0_6_33;   // mult_24u_24u.v(405[10:31])
    wire s_mult_24u_24u_0_7_34;   // mult_24u_24u.v(404[10:31])
    wire s_mult_24u_24u_0_7_33;   // mult_24u_24u.v(403[10:31])
    wire co_mult_24u_24u_0_9_13;   // mult_24u_24u.v(402[10:32])
    wire s_mult_24u_24u_0_6_32;   // mult_24u_24u.v(401[10:31])
    wire s_mult_24u_24u_0_6_31;   // mult_24u_24u.v(400[10:31])
    wire s_mult_24u_24u_0_7_32;   // mult_24u_24u.v(399[10:31])
    wire s_mult_24u_24u_0_7_31;   // mult_24u_24u.v(398[10:31])
    wire co_mult_24u_24u_0_9_12;   // mult_24u_24u.v(397[10:32])
    wire s_mult_24u_24u_0_6_30;   // mult_24u_24u.v(396[10:31])
    wire s_mult_24u_24u_0_6_29;   // mult_24u_24u.v(395[10:31])
    wire s_mult_24u_24u_0_7_30;   // mult_24u_24u.v(394[10:31])
    wire s_mult_24u_24u_0_7_29;   // mult_24u_24u.v(393[10:31])
    wire co_mult_24u_24u_0_9_11;   // mult_24u_24u.v(392[10:32])
    wire s_mult_24u_24u_0_6_28;   // mult_24u_24u.v(391[10:31])
    wire s_mult_24u_24u_0_6_27;   // mult_24u_24u.v(390[10:31])
    wire s_mult_24u_24u_0_7_28;   // mult_24u_24u.v(389[10:31])
    wire s_mult_24u_24u_0_7_27;   // mult_24u_24u.v(388[10:31])
    wire co_mult_24u_24u_0_9_10;   // mult_24u_24u.v(387[10:32])
    wire s_mult_24u_24u_0_6_26;   // mult_24u_24u.v(386[10:31])
    wire s_mult_24u_24u_0_6_25;   // mult_24u_24u.v(385[10:31])
    wire s_mult_24u_24u_0_7_26;   // mult_24u_24u.v(384[10:31])
    wire s_mult_24u_24u_0_7_25;   // mult_24u_24u.v(383[10:31])
    wire co_mult_24u_24u_0_9_9;   // mult_24u_24u.v(382[10:31])
    wire s_mult_24u_24u_0_6_24;   // mult_24u_24u.v(381[10:31])
    wire s_mult_24u_24u_0_6_23;   // mult_24u_24u.v(380[10:31])
    wire s_mult_24u_24u_0_7_24;   // mult_24u_24u.v(379[10:31])
    wire s_mult_24u_24u_0_7_23;   // mult_24u_24u.v(378[10:31])
    wire co_mult_24u_24u_0_9_8;   // mult_24u_24u.v(377[10:31])
    wire s_mult_24u_24u_0_6_22;   // mult_24u_24u.v(376[10:31])
    wire s_mult_24u_24u_0_6_21;   // mult_24u_24u.v(375[10:31])
    wire s_mult_24u_24u_0_7_22;   // mult_24u_24u.v(374[10:31])
    wire s_mult_24u_24u_0_7_21;   // mult_24u_24u.v(373[10:31])
    wire co_mult_24u_24u_0_9_7;   // mult_24u_24u.v(372[10:31])
    wire s_mult_24u_24u_0_6_20;   // mult_24u_24u.v(371[10:31])
    wire s_mult_24u_24u_0_6_19;   // mult_24u_24u.v(370[10:31])
    wire s_mult_24u_24u_0_7_20;   // mult_24u_24u.v(369[10:31])
    wire s_mult_24u_24u_0_7_19;   // mult_24u_24u.v(368[10:31])
    wire co_mult_24u_24u_0_9_6;   // mult_24u_24u.v(367[10:31])
    wire s_mult_24u_24u_0_6_18;   // mult_24u_24u.v(366[10:31])
    wire s_mult_24u_24u_0_6_17;   // mult_24u_24u.v(365[10:31])
    wire s_mult_24u_24u_0_7_18;   // mult_24u_24u.v(364[10:31])
    wire s_mult_24u_24u_0_7_17;   // mult_24u_24u.v(363[10:31])
    wire co_mult_24u_24u_0_9_5;   // mult_24u_24u.v(362[10:31])
    wire s_mult_24u_24u_0_6_16;   // mult_24u_24u.v(361[10:31])
    wire s_mult_24u_24u_0_6_15;   // mult_24u_24u.v(360[10:31])
    wire s_mult_24u_24u_0_7_16;   // mult_24u_24u.v(359[10:31])
    wire s_mult_24u_24u_0_7_15;   // mult_24u_24u.v(358[10:31])
    wire co_mult_24u_24u_0_9_4;   // mult_24u_24u.v(357[10:31])
    wire s_mult_24u_24u_0_6_14;   // mult_24u_24u.v(355[10:31])
    wire s_mult_24u_24u_0_6_13;   // mult_24u_24u.v(354[10:31])
    wire s_mult_24u_24u_0_7_14;   // mult_24u_24u.v(353[10:31])
    wire s_mult_24u_24u_0_7_13;   // mult_24u_24u.v(352[10:31])
    wire co_mult_24u_24u_0_9_3;   // mult_24u_24u.v(351[10:31])
    wire s_mult_24u_24u_0_6_12;   // mult_24u_24u.v(348[10:31])
    wire s_mult_24u_24u_0_6_11;   // mult_24u_24u.v(347[10:31])
    wire s_mult_24u_24u_0_7_12;   // mult_24u_24u.v(346[10:31])
    wire s_mult_24u_24u_0_2_11;   // mult_24u_24u.v(345[10:31])
    wire co_mult_24u_24u_0_9_2;   // mult_24u_24u.v(344[10:31])
    wire s_mult_24u_24u_0_6_10;   // mult_24u_24u.v(341[10:31])
    wire s_mult_24u_24u_0_6_9;   // mult_24u_24u.v(340[10:30])
    wire s_mult_24u_24u_0_2_10;   // mult_24u_24u.v(339[10:31])
    wire co_mult_24u_24u_0_9_1;   // mult_24u_24u.v(338[10:31])
    wire s_mult_24u_24u_0_6_8;   // mult_24u_24u.v(335[10:30])
    wire mult_24u_24u_0_pp_4_8;   // mult_24u_24u.v(334[10:31])
    wire s_mult_24u_24u_0_5_47;   // mult_24u_24u.v(332[10:31])
    wire co_mult_24u_24u_0_8_14;   // mult_24u_24u.v(331[10:32])
    wire s_mult_24u_24u_0_4_45;   // mult_24u_24u.v(329[10:31])
    wire s_mult_24u_24u_0_5_46;   // mult_24u_24u.v(328[10:31])
    wire s_mult_24u_24u_0_5_45;   // mult_24u_24u.v(327[10:31])
    wire co_mult_24u_24u_0_8_13;   // mult_24u_24u.v(326[10:32])
    wire s_mult_24u_24u_0_4_44;   // mult_24u_24u.v(325[10:31])
    wire s_mult_24u_24u_0_4_43;   // mult_24u_24u.v(324[10:31])
    wire s_mult_24u_24u_0_5_44;   // mult_24u_24u.v(323[10:31])
    wire s_mult_24u_24u_0_5_43;   // mult_24u_24u.v(322[10:31])
    wire co_mult_24u_24u_0_8_12;   // mult_24u_24u.v(321[10:32])
    wire s_mult_24u_24u_0_4_42;   // mult_24u_24u.v(320[10:31])
    wire s_mult_24u_24u_0_4_41;   // mult_24u_24u.v(319[10:31])
    wire s_mult_24u_24u_0_5_42;   // mult_24u_24u.v(318[10:31])
    wire s_mult_24u_24u_0_5_41;   // mult_24u_24u.v(317[10:31])
    wire co_mult_24u_24u_0_8_11;   // mult_24u_24u.v(316[10:32])
    wire s_mult_24u_24u_0_4_40;   // mult_24u_24u.v(315[10:31])
    wire s_mult_24u_24u_0_4_39;   // mult_24u_24u.v(314[10:31])
    wire s_mult_24u_24u_0_5_40;   // mult_24u_24u.v(313[10:31])
    wire s_mult_24u_24u_0_5_39;   // mult_24u_24u.v(312[10:31])
    wire co_mult_24u_24u_0_8_10;   // mult_24u_24u.v(311[10:32])
    wire s_mult_24u_24u_0_4_38;   // mult_24u_24u.v(310[10:31])
    wire s_mult_24u_24u_0_4_37;   // mult_24u_24u.v(309[10:31])
    wire s_mult_24u_24u_0_5_38;   // mult_24u_24u.v(308[10:31])
    wire s_mult_24u_24u_0_5_37;   // mult_24u_24u.v(307[10:31])
    wire co_mult_24u_24u_0_8_9;   // mult_24u_24u.v(306[10:31])
    wire s_mult_24u_24u_0_4_36;   // mult_24u_24u.v(305[10:31])
    wire s_mult_24u_24u_0_4_35;   // mult_24u_24u.v(304[10:31])
    wire s_mult_24u_24u_0_5_36;   // mult_24u_24u.v(303[10:31])
    wire s_mult_24u_24u_0_5_35;   // mult_24u_24u.v(302[10:31])
    wire co_mult_24u_24u_0_8_8;   // mult_24u_24u.v(301[10:31])
    wire s_mult_24u_24u_0_4_34;   // mult_24u_24u.v(300[10:31])
    wire s_mult_24u_24u_0_4_33;   // mult_24u_24u.v(299[10:31])
    wire s_mult_24u_24u_0_5_34;   // mult_24u_24u.v(298[10:31])
    wire s_mult_24u_24u_0_5_33;   // mult_24u_24u.v(297[10:31])
    wire co_mult_24u_24u_0_8_7;   // mult_24u_24u.v(296[10:31])
    wire s_mult_24u_24u_0_4_32;   // mult_24u_24u.v(295[10:31])
    wire s_mult_24u_24u_0_4_31;   // mult_24u_24u.v(294[10:31])
    wire s_mult_24u_24u_0_5_32;   // mult_24u_24u.v(293[10:31])
    wire s_mult_24u_24u_0_5_31;   // mult_24u_24u.v(292[10:31])
    wire co_mult_24u_24u_0_8_6;   // mult_24u_24u.v(291[10:31])
    wire s_mult_24u_24u_0_4_30;   // mult_24u_24u.v(290[10:31])
    wire s_mult_24u_24u_0_4_29;   // mult_24u_24u.v(289[10:31])
    wire s_mult_24u_24u_0_5_30;   // mult_24u_24u.v(288[10:31])
    wire s_mult_24u_24u_0_5_29;   // mult_24u_24u.v(287[10:31])
    wire co_mult_24u_24u_0_8_5;   // mult_24u_24u.v(286[10:31])
    wire s_mult_24u_24u_0_4_28;   // mult_24u_24u.v(285[10:31])
    wire s_mult_24u_24u_0_4_27;   // mult_24u_24u.v(284[10:31])
    wire s_mult_24u_24u_0_5_28;   // mult_24u_24u.v(283[10:31])
    wire s_mult_24u_24u_0_5_27;   // mult_24u_24u.v(282[10:31])
    wire co_mult_24u_24u_0_8_4;   // mult_24u_24u.v(281[10:31])
    wire s_mult_24u_24u_0_4_26;   // mult_24u_24u.v(280[10:31])
    wire s_mult_24u_24u_0_4_25;   // mult_24u_24u.v(279[10:31])
    wire s_mult_24u_24u_0_5_26;   // mult_24u_24u.v(278[10:31])
    wire s_mult_24u_24u_0_5_25;   // mult_24u_24u.v(277[10:31])
    wire co_mult_24u_24u_0_8_3;   // mult_24u_24u.v(276[10:31])
    wire s_mult_24u_24u_0_4_24;   // mult_24u_24u.v(275[10:31])
    wire s_mult_24u_24u_0_4_23;   // mult_24u_24u.v(274[10:31])
    wire s_mult_24u_24u_0_5_24;   // mult_24u_24u.v(273[10:31])
    wire s_mult_24u_24u_0_5_23;   // mult_24u_24u.v(272[10:31])
    wire co_mult_24u_24u_0_8_2;   // mult_24u_24u.v(271[10:31])
    wire s_mult_24u_24u_0_4_22;   // mult_24u_24u.v(270[10:31])
    wire s_mult_24u_24u_0_4_21;   // mult_24u_24u.v(269[10:31])
    wire s_mult_24u_24u_0_5_22;   // mult_24u_24u.v(268[10:31])
    wire co_mult_24u_24u_0_8_1;   // mult_24u_24u.v(267[10:31])
    wire s_mult_24u_24u_0_4_20;   // mult_24u_24u.v(266[10:31])
    wire mult_24u_24u_0_pp_10_20;   // mult_24u_24u.v(265[10:33])
    wire co_mult_24u_24u_0_7_16;   // mult_24u_24u.v(264[10:32])
    wire s_mult_24u_24u_0_3_41;   // mult_24u_24u.v(263[10:31])
    wire co_mult_24u_24u_0_7_15;   // mult_24u_24u.v(262[10:32])
    wire s_mult_24u_24u_0_3_40;   // mult_24u_24u.v(261[10:31])
    wire s_mult_24u_24u_0_3_39;   // mult_24u_24u.v(260[10:31])
    wire co_mult_24u_24u_0_7_14;   // mult_24u_24u.v(259[10:32])
    wire s_mult_24u_24u_0_2_37;   // mult_24u_24u.v(258[10:31])
    wire s_mult_24u_24u_0_3_38;   // mult_24u_24u.v(257[10:31])
    wire s_mult_24u_24u_0_3_37;   // mult_24u_24u.v(256[10:31])
    wire co_mult_24u_24u_0_7_13;   // mult_24u_24u.v(255[10:32])
    wire s_mult_24u_24u_0_2_36;   // mult_24u_24u.v(254[10:31])
    wire s_mult_24u_24u_0_2_35;   // mult_24u_24u.v(253[10:31])
    wire s_mult_24u_24u_0_3_36;   // mult_24u_24u.v(252[10:31])
    wire s_mult_24u_24u_0_3_35;   // mult_24u_24u.v(251[10:31])
    wire co_mult_24u_24u_0_7_12;   // mult_24u_24u.v(250[10:32])
    wire s_mult_24u_24u_0_2_34;   // mult_24u_24u.v(249[10:31])
    wire s_mult_24u_24u_0_2_33;   // mult_24u_24u.v(248[10:31])
    wire s_mult_24u_24u_0_3_34;   // mult_24u_24u.v(247[10:31])
    wire s_mult_24u_24u_0_3_33;   // mult_24u_24u.v(246[10:31])
    wire co_mult_24u_24u_0_7_11;   // mult_24u_24u.v(245[10:32])
    wire s_mult_24u_24u_0_2_32;   // mult_24u_24u.v(244[10:31])
    wire s_mult_24u_24u_0_2_31;   // mult_24u_24u.v(243[10:31])
    wire s_mult_24u_24u_0_3_32;   // mult_24u_24u.v(242[10:31])
    wire s_mult_24u_24u_0_3_31;   // mult_24u_24u.v(241[10:31])
    wire co_mult_24u_24u_0_7_10;   // mult_24u_24u.v(240[10:32])
    wire s_mult_24u_24u_0_2_30;   // mult_24u_24u.v(239[10:31])
    wire s_mult_24u_24u_0_2_29;   // mult_24u_24u.v(238[10:31])
    wire s_mult_24u_24u_0_3_30;   // mult_24u_24u.v(237[10:31])
    wire s_mult_24u_24u_0_3_29;   // mult_24u_24u.v(236[10:31])
    wire co_mult_24u_24u_0_7_9;   // mult_24u_24u.v(235[10:31])
    wire s_mult_24u_24u_0_2_28;   // mult_24u_24u.v(234[10:31])
    wire s_mult_24u_24u_0_2_27;   // mult_24u_24u.v(233[10:31])
    wire s_mult_24u_24u_0_3_28;   // mult_24u_24u.v(232[10:31])
    wire s_mult_24u_24u_0_3_27;   // mult_24u_24u.v(231[10:31])
    wire co_mult_24u_24u_0_7_8;   // mult_24u_24u.v(230[10:31])
    wire s_mult_24u_24u_0_2_26;   // mult_24u_24u.v(229[10:31])
    wire s_mult_24u_24u_0_2_25;   // mult_24u_24u.v(228[10:31])
    wire s_mult_24u_24u_0_3_26;   // mult_24u_24u.v(227[10:31])
    wire s_mult_24u_24u_0_3_25;   // mult_24u_24u.v(226[10:31])
    wire co_mult_24u_24u_0_7_7;   // mult_24u_24u.v(225[10:31])
    wire s_mult_24u_24u_0_2_24;   // mult_24u_24u.v(224[10:31])
    wire s_mult_24u_24u_0_2_23;   // mult_24u_24u.v(223[10:31])
    wire s_mult_24u_24u_0_3_24;   // mult_24u_24u.v(222[10:31])
    wire s_mult_24u_24u_0_3_23;   // mult_24u_24u.v(221[10:31])
    wire co_mult_24u_24u_0_7_6;   // mult_24u_24u.v(220[10:31])
    wire s_mult_24u_24u_0_2_22;   // mult_24u_24u.v(219[10:31])
    wire s_mult_24u_24u_0_2_21;   // mult_24u_24u.v(218[10:31])
    wire s_mult_24u_24u_0_3_22;   // mult_24u_24u.v(217[10:31])
    wire s_mult_24u_24u_0_3_21;   // mult_24u_24u.v(216[10:31])
    wire co_mult_24u_24u_0_7_5;   // mult_24u_24u.v(215[10:31])
    wire s_mult_24u_24u_0_2_20;   // mult_24u_24u.v(214[10:31])
    wire s_mult_24u_24u_0_2_19;   // mult_24u_24u.v(213[10:31])
    wire s_mult_24u_24u_0_3_20;   // mult_24u_24u.v(212[10:31])
    wire s_mult_24u_24u_0_3_19;   // mult_24u_24u.v(211[10:31])
    wire co_mult_24u_24u_0_7_4;   // mult_24u_24u.v(210[10:31])
    wire s_mult_24u_24u_0_2_18;   // mult_24u_24u.v(209[10:31])
    wire s_mult_24u_24u_0_2_17;   // mult_24u_24u.v(208[10:31])
    wire s_mult_24u_24u_0_3_18;   // mult_24u_24u.v(207[10:31])
    wire s_mult_24u_24u_0_3_17;   // mult_24u_24u.v(206[10:31])
    wire co_mult_24u_24u_0_7_3;   // mult_24u_24u.v(205[10:31])
    wire s_mult_24u_24u_0_2_16;   // mult_24u_24u.v(204[10:31])
    wire s_mult_24u_24u_0_2_15;   // mult_24u_24u.v(203[10:31])
    wire s_mult_24u_24u_0_3_16;   // mult_24u_24u.v(202[10:31])
    wire s_mult_24u_24u_0_3_15;   // mult_24u_24u.v(201[10:31])
    wire co_mult_24u_24u_0_7_2;   // mult_24u_24u.v(200[10:31])
    wire s_mult_24u_24u_0_2_14;   // mult_24u_24u.v(199[10:31])
    wire s_mult_24u_24u_0_2_13;   // mult_24u_24u.v(198[10:31])
    wire s_mult_24u_24u_0_3_14;   // mult_24u_24u.v(197[10:31])
    wire co_mult_24u_24u_0_7_1;   // mult_24u_24u.v(196[10:31])
    wire s_mult_24u_24u_0_2_12;   // mult_24u_24u.v(195[10:31])
    wire mult_24u_24u_0_pp_6_12;   // mult_24u_24u.v(194[10:32])
    wire co_mult_24u_24u_0_6_16;   // mult_24u_24u.v(193[10:32])
    wire s_mult_24u_24u_0_1_33;   // mult_24u_24u.v(192[10:31])
    wire co_mult_24u_24u_0_6_15;   // mult_24u_24u.v(191[10:32])
    wire s_mult_24u_24u_0_1_32;   // mult_24u_24u.v(190[10:31])
    wire s_mult_24u_24u_0_1_31;   // mult_24u_24u.v(189[10:31])
    wire co_mult_24u_24u_0_6_14;   // mult_24u_24u.v(188[10:32])
    wire s_mult_24u_24u_0_0_29;   // mult_24u_24u.v(187[10:31])
    wire s_mult_24u_24u_0_1_30;   // mult_24u_24u.v(186[10:31])
    wire s_mult_24u_24u_0_1_29;   // mult_24u_24u.v(185[10:31])
    wire co_mult_24u_24u_0_6_13;   // mult_24u_24u.v(184[10:32])
    wire s_mult_24u_24u_0_0_28;   // mult_24u_24u.v(183[10:31])
    wire s_mult_24u_24u_0_0_27;   // mult_24u_24u.v(182[10:31])
    wire s_mult_24u_24u_0_1_28;   // mult_24u_24u.v(181[10:31])
    wire s_mult_24u_24u_0_1_27;   // mult_24u_24u.v(180[10:31])
    wire co_mult_24u_24u_0_6_12;   // mult_24u_24u.v(179[10:32])
    wire s_mult_24u_24u_0_0_26;   // mult_24u_24u.v(178[10:31])
    wire s_mult_24u_24u_0_0_25;   // mult_24u_24u.v(177[10:31])
    wire s_mult_24u_24u_0_1_26;   // mult_24u_24u.v(176[10:31])
    wire s_mult_24u_24u_0_1_25;   // mult_24u_24u.v(175[10:31])
    wire co_mult_24u_24u_0_6_11;   // mult_24u_24u.v(174[10:32])
    wire s_mult_24u_24u_0_0_24;   // mult_24u_24u.v(173[10:31])
    wire s_mult_24u_24u_0_0_23;   // mult_24u_24u.v(172[10:31])
    wire s_mult_24u_24u_0_1_24;   // mult_24u_24u.v(171[10:31])
    wire s_mult_24u_24u_0_1_23;   // mult_24u_24u.v(170[10:31])
    wire co_mult_24u_24u_0_6_10;   // mult_24u_24u.v(169[10:32])
    wire s_mult_24u_24u_0_0_22;   // mult_24u_24u.v(168[10:31])
    wire s_mult_24u_24u_0_0_21;   // mult_24u_24u.v(167[10:31])
    wire s_mult_24u_24u_0_1_22;   // mult_24u_24u.v(166[10:31])
    wire s_mult_24u_24u_0_1_21;   // mult_24u_24u.v(165[10:31])
    wire co_mult_24u_24u_0_6_9;   // mult_24u_24u.v(164[10:31])
    wire s_mult_24u_24u_0_0_20;   // mult_24u_24u.v(163[10:31])
    wire s_mult_24u_24u_0_0_19;   // mult_24u_24u.v(162[10:31])
    wire s_mult_24u_24u_0_1_20;   // mult_24u_24u.v(161[10:31])
    wire s_mult_24u_24u_0_1_19;   // mult_24u_24u.v(160[10:31])
    wire co_mult_24u_24u_0_6_8;   // mult_24u_24u.v(159[10:31])
    wire s_mult_24u_24u_0_0_18;   // mult_24u_24u.v(158[10:31])
    wire s_mult_24u_24u_0_0_17;   // mult_24u_24u.v(157[10:31])
    wire s_mult_24u_24u_0_1_18;   // mult_24u_24u.v(156[10:31])
    wire s_mult_24u_24u_0_1_17;   // mult_24u_24u.v(155[10:31])
    wire co_mult_24u_24u_0_6_7;   // mult_24u_24u.v(154[10:31])
    wire s_mult_24u_24u_0_0_16;   // mult_24u_24u.v(153[10:31])
    wire s_mult_24u_24u_0_0_15;   // mult_24u_24u.v(152[10:31])
    wire s_mult_24u_24u_0_1_16;   // mult_24u_24u.v(151[10:31])
    wire s_mult_24u_24u_0_1_15;   // mult_24u_24u.v(150[10:31])
    wire co_mult_24u_24u_0_6_6;   // mult_24u_24u.v(149[10:31])
    wire s_mult_24u_24u_0_0_14;   // mult_24u_24u.v(148[10:31])
    wire s_mult_24u_24u_0_0_13;   // mult_24u_24u.v(147[10:31])
    wire s_mult_24u_24u_0_1_14;   // mult_24u_24u.v(146[10:31])
    wire s_mult_24u_24u_0_1_13;   // mult_24u_24u.v(145[10:31])
    wire co_mult_24u_24u_0_6_5;   // mult_24u_24u.v(144[10:31])
    wire s_mult_24u_24u_0_0_12;   // mult_24u_24u.v(143[10:31])
    wire s_mult_24u_24u_0_0_11;   // mult_24u_24u.v(142[10:31])
    wire s_mult_24u_24u_0_1_12;   // mult_24u_24u.v(141[10:31])
    wire s_mult_24u_24u_0_1_11;   // mult_24u_24u.v(140[10:31])
    wire co_mult_24u_24u_0_6_4;   // mult_24u_24u.v(139[10:31])
    wire s_mult_24u_24u_0_0_10;   // mult_24u_24u.v(138[10:31])
    wire s_mult_24u_24u_0_0_9;   // mult_24u_24u.v(137[10:30])
    wire s_mult_24u_24u_0_1_10;   // mult_24u_24u.v(136[10:31])
    wire s_mult_24u_24u_0_1_9;   // mult_24u_24u.v(135[10:30])
    wire co_mult_24u_24u_0_6_3;   // mult_24u_24u.v(134[10:31])
    wire s_mult_24u_24u_0_0_8;   // mult_24u_24u.v(133[10:30])
    wire s_mult_24u_24u_0_0_7;   // mult_24u_24u.v(132[10:30])
    wire s_mult_24u_24u_0_1_8;   // mult_24u_24u.v(131[10:30])
    wire s_mult_24u_24u_0_1_7;   // mult_24u_24u.v(130[10:30])
    wire co_mult_24u_24u_0_6_2;   // mult_24u_24u.v(129[10:31])
    wire s_mult_24u_24u_0_0_6;   // mult_24u_24u.v(127[10:30])
    wire s_mult_24u_24u_0_0_5;   // mult_24u_24u.v(126[10:30])
    wire s_mult_24u_24u_0_1_6;   // mult_24u_24u.v(125[10:30])
    wire co_mult_24u_24u_0_6_1;   // mult_24u_24u.v(124[10:31])
    wire s_mult_24u_24u_0_0_4;   // mult_24u_24u.v(121[10:30])
    wire mult_24u_24u_0_pp_2_4;   // mult_24u_24u.v(120[10:31])
    wire mult_24u_24u_0_pp_11_47;   // mult_24u_24u.v(118[10:33])
    wire co_mult_24u_24u_0_5_13;   // mult_24u_24u.v(117[10:32])
    wire mult_24u_24u_0_pp_10_45;   // mult_24u_24u.v(115[10:33])
    wire co_mult_24u_24u_0_5_12;   // mult_24u_24u.v(114[10:32])
    wire co_mult_24u_24u_0_5_11;   // mult_24u_24u.v(113[10:32])
    wire co_mult_24u_24u_0_5_10;   // mult_24u_24u.v(112[10:32])
    wire co_mult_24u_24u_0_5_9;   // mult_24u_24u.v(111[10:31])
    wire co_mult_24u_24u_0_5_8;   // mult_24u_24u.v(110[10:31])
    wire co_mult_24u_24u_0_5_7;   // mult_24u_24u.v(109[10:31])
    wire co_mult_24u_24u_0_5_6;   // mult_24u_24u.v(108[10:31])
    wire co_mult_24u_24u_0_5_5;   // mult_24u_24u.v(107[10:31])
    wire co_mult_24u_24u_0_5_4;   // mult_24u_24u.v(106[10:31])
    wire co_mult_24u_24u_0_5_3;   // mult_24u_24u.v(105[10:31])
    wire co_mult_24u_24u_0_5_2;   // mult_24u_24u.v(104[10:31])
    wire co_mult_24u_24u_0_5_1;   // mult_24u_24u.v(103[10:31])
    wire mult_24u_24u_0_pp_11_22;   // mult_24u_24u.v(102[10:33])
    wire co_mult_24u_24u_0_4_14;   // mult_24u_24u.v(101[10:32])
    wire mult_24u_24u_0_pp_9_43;   // mult_24u_24u.v(100[10:32])
    wire co_mult_24u_24u_0_4_13;   // mult_24u_24u.v(99[10:32])
    wire mult_24u_24u_0_pp_8_41;   // mult_24u_24u.v(98[10:32])
    wire co_mult_24u_24u_0_4_12;   // mult_24u_24u.v(97[10:32])
    wire co_mult_24u_24u_0_4_11;   // mult_24u_24u.v(96[10:32])
    wire co_mult_24u_24u_0_4_10;   // mult_24u_24u.v(95[10:32])
    wire co_mult_24u_24u_0_4_9;   // mult_24u_24u.v(94[10:31])
    wire co_mult_24u_24u_0_4_8;   // mult_24u_24u.v(93[10:31])
    wire co_mult_24u_24u_0_4_7;   // mult_24u_24u.v(92[10:31])
    wire co_mult_24u_24u_0_4_6;   // mult_24u_24u.v(91[10:31])
    wire co_mult_24u_24u_0_4_5;   // mult_24u_24u.v(90[10:31])
    wire co_mult_24u_24u_0_4_4;   // mult_24u_24u.v(89[10:31])
    wire co_mult_24u_24u_0_4_3;   // mult_24u_24u.v(88[10:31])
    wire co_mult_24u_24u_0_4_2;   // mult_24u_24u.v(87[10:31])
    wire co_mult_24u_24u_0_4_1;   // mult_24u_24u.v(86[10:31])
    wire mult_24u_24u_0_pp_9_18;   // mult_24u_24u.v(85[10:32])
    wire co_mult_24u_24u_0_3_14;   // mult_24u_24u.v(84[10:32])
    wire mult_24u_24u_0_pp_7_39;   // mult_24u_24u.v(83[10:32])
    wire co_mult_24u_24u_0_3_13;   // mult_24u_24u.v(82[10:32])
    wire mult_24u_24u_0_pp_6_37;   // mult_24u_24u.v(81[10:32])
    wire co_mult_24u_24u_0_3_12;   // mult_24u_24u.v(80[10:32])
    wire co_mult_24u_24u_0_3_11;   // mult_24u_24u.v(79[10:32])
    wire co_mult_24u_24u_0_3_10;   // mult_24u_24u.v(78[10:32])
    wire co_mult_24u_24u_0_3_9;   // mult_24u_24u.v(77[10:31])
    wire co_mult_24u_24u_0_3_8;   // mult_24u_24u.v(76[10:31])
    wire co_mult_24u_24u_0_3_7;   // mult_24u_24u.v(75[10:31])
    wire co_mult_24u_24u_0_3_6;   // mult_24u_24u.v(74[10:31])
    wire co_mult_24u_24u_0_3_5;   // mult_24u_24u.v(73[10:31])
    wire co_mult_24u_24u_0_3_4;   // mult_24u_24u.v(72[10:31])
    wire co_mult_24u_24u_0_3_3;   // mult_24u_24u.v(71[10:31])
    wire co_mult_24u_24u_0_3_2;   // mult_24u_24u.v(70[10:31])
    wire co_mult_24u_24u_0_3_1;   // mult_24u_24u.v(69[10:31])
    wire mult_24u_24u_0_pp_7_14;   // mult_24u_24u.v(68[10:32])
    wire co_mult_24u_24u_0_2_14;   // mult_24u_24u.v(67[10:32])
    wire mult_24u_24u_0_pp_5_35;   // mult_24u_24u.v(66[10:32])
    wire co_mult_24u_24u_0_2_13;   // mult_24u_24u.v(65[10:32])
    wire mult_24u_24u_0_pp_4_33;   // mult_24u_24u.v(64[10:32])
    wire co_mult_24u_24u_0_2_12;   // mult_24u_24u.v(63[10:32])
    wire co_mult_24u_24u_0_2_11;   // mult_24u_24u.v(62[10:32])
    wire co_mult_24u_24u_0_2_10;   // mult_24u_24u.v(61[10:32])
    wire co_mult_24u_24u_0_2_9;   // mult_24u_24u.v(60[10:31])
    wire co_mult_24u_24u_0_2_8;   // mult_24u_24u.v(59[10:31])
    wire co_mult_24u_24u_0_2_7;   // mult_24u_24u.v(58[10:31])
    wire co_mult_24u_24u_0_2_6;   // mult_24u_24u.v(57[10:31])
    wire co_mult_24u_24u_0_2_5;   // mult_24u_24u.v(56[10:31])
    wire co_mult_24u_24u_0_2_4;   // mult_24u_24u.v(55[10:31])
    wire co_mult_24u_24u_0_2_3;   // mult_24u_24u.v(54[10:31])
    wire co_mult_24u_24u_0_2_2;   // mult_24u_24u.v(53[10:31])
    wire co_mult_24u_24u_0_2_1;   // mult_24u_24u.v(52[10:31])
    wire mult_24u_24u_0_pp_5_10;   // mult_24u_24u.v(51[10:32])
    wire co_mult_24u_24u_0_1_14;   // mult_24u_24u.v(50[10:32])
    wire mult_24u_24u_0_pp_3_31;   // mult_24u_24u.v(49[10:32])
    wire co_mult_24u_24u_0_1_13;   // mult_24u_24u.v(48[10:32])
    wire mult_24u_24u_0_pp_2_29;   // mult_24u_24u.v(47[10:32])
    wire co_mult_24u_24u_0_1_12;   // mult_24u_24u.v(46[10:32])
    wire co_mult_24u_24u_0_1_11;   // mult_24u_24u.v(45[10:32])
    wire co_mult_24u_24u_0_1_10;   // mult_24u_24u.v(44[10:32])
    wire co_mult_24u_24u_0_1_9;   // mult_24u_24u.v(43[10:31])
    wire co_mult_24u_24u_0_1_8;   // mult_24u_24u.v(42[10:31])
    wire co_mult_24u_24u_0_1_7;   // mult_24u_24u.v(41[10:31])
    wire co_mult_24u_24u_0_1_6;   // mult_24u_24u.v(40[10:31])
    wire co_mult_24u_24u_0_1_5;   // mult_24u_24u.v(39[10:31])
    wire co_mult_24u_24u_0_1_4;   // mult_24u_24u.v(38[10:31])
    wire co_mult_24u_24u_0_1_3;   // mult_24u_24u.v(37[10:31])
    wire co_mult_24u_24u_0_1_2;   // mult_24u_24u.v(36[10:31])
    wire co_mult_24u_24u_0_1_1;   // mult_24u_24u.v(35[10:31])
    wire mult_24u_24u_0_pp_3_6;   // mult_24u_24u.v(34[10:31])
    wire co_mult_24u_24u_0_0_14;   // mult_24u_24u.v(33[10:32])
    wire mult_24u_24u_0_pp_1_27;   // mult_24u_24u.v(32[10:32])
    wire co_mult_24u_24u_0_0_13;   // mult_24u_24u.v(31[10:32])
    wire mult_24u_24u_0_pp_0_25;   // mult_24u_24u.v(30[10:32])
    wire co_mult_24u_24u_0_0_12;   // mult_24u_24u.v(29[10:32])
    wire co_mult_24u_24u_0_0_11;   // mult_24u_24u.v(28[10:32])
    wire co_mult_24u_24u_0_0_10;   // mult_24u_24u.v(27[10:32])
    wire co_mult_24u_24u_0_0_9;   // mult_24u_24u.v(26[10:31])
    wire co_mult_24u_24u_0_0_8;   // mult_24u_24u.v(25[10:31])
    wire co_mult_24u_24u_0_0_7;   // mult_24u_24u.v(24[10:31])
    wire co_mult_24u_24u_0_0_6;   // mult_24u_24u.v(23[10:31])
    wire co_mult_24u_24u_0_0_5;   // mult_24u_24u.v(22[10:31])
    wire co_mult_24u_24u_0_0_4;   // mult_24u_24u.v(21[10:31])
    wire co_mult_24u_24u_0_0_3;   // mult_24u_24u.v(20[10:31])
    wire co_mult_24u_24u_0_0_2;   // mult_24u_24u.v(19[10:31])
    wire co_mult_24u_24u_0_0_1;   // mult_24u_24u.v(18[10:31])
    wire mult_24u_24u_0_pp_1_2;   // mult_24u_24u.v(16[10:31])
    wire mco_adj_571;   // mult_2u_3u.v(21[10:13])
    wire mult_2u_3u_0_cin_lr_0;   // mult_2u_3u.v(17[10:31])
    wire mco_adj_572;   // mult_3u_2u.v(21[10:13])
    wire mult_3u_2u_0_cin_lr_0;   // mult_3u_2u.v(17[10:31])
    wire mult_2u_2u_0_cin_lr_0;   // mult_2u_2u.v(19[10:31])
    wire mfco_adj_573;   // mult_2u_2u.v(16[10:14])
    wire [1:0]state_adj_642;   // c:/users/yisong/documents/new/mlp/pr.vhd(30[8:13])
    wire spi_mosi_oe;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(35[12:23])
    wire spi_mosi_o;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(36[12:22])
    wire spi_miso_oe;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(37[12:23])
    wire spi_miso_o;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(38[12:22])
    wire spi_clk_oe;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(39[12:22])
    wire spi_clk_o;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(40[12:21])
    wire spi_mosi_i;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(41[12:22])
    wire spi_miso_i;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(42[12:22])
    wire spi_clk_i;   // c:/users/yisong/documents/new/mlp/efb_spi.vhd(43[12:21])
    wire [31:0]A_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(54[11:16])
    wire [31:0]B_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(55[11:16])
    wire [27:0]efectFracB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(67[23:33])
    wire [8:0]diffExpAB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[11:20])
    wire [8:0]diffExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[33:40])
    wire [31:0]A_int_adj_660;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(54[11:16])
    wire [31:0]B_int_adj_661;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(55[11:16])
    wire [27:0]efectFracB_adj_666;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(67[23:33])
    wire [8:0]diffExpAB_adj_668;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[11:20])
    wire [27:0]frac_adj_677;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(97[11:15])
    wire [31:0]A_int_adj_724;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(44[11:16])
    wire [31:0]B_int_adj_725;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(44[18:23])
    wire [47:0]prod;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(53[11:15])
    wire [26:0]frac_norm;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(63[11:20])
    wire [7:0]exp_final;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(68[11:20])
    wire [31:0]FP_Z_int_adj_729;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(69[11:19])
    wire [1:0]n14053;   // mult_2u_3u.v(10[22:23])
    wire [33:0]n898;   // mult_32s_2s.v(11[24:25])
    wire [166:0]buf_x_adj_1109;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [166:0]buf_r_adj_1110;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(337[10:15])
    wire [1:0]n14049;   // mult_3u_2u.v(9[22:23])
    wire n73802 /* synthesis nomerge= */ ;
    wire mult_32s_2s_0_cin_lr;   // mult_32s_2s.v(18[10:30])
    wire mult_32s_2s_0_mult_0_0_n1;   // mult_32s_2s.v(19[10:35])
    wire mult_32s_2s_0_mult_0_0_n0;   // mult_32s_2s.v(20[10:35])
    wire mco_adj_608;   // mult_32s_2s.v(23[10:13])
    wire mult_32s_2s_0_mult_0_1_n1;   // mult_32s_2s.v(24[10:35])
    wire mult_32s_2s_0_mult_0_1_n0;   // mult_32s_2s.v(25[10:35])
    wire mco_1_adj_609;   // mult_32s_2s.v(28[10:15])
    wire mult_32s_2s_0_mult_0_2_n1;   // mult_32s_2s.v(29[10:35])
    wire mult_32s_2s_0_mult_0_2_n0;   // mult_32s_2s.v(30[10:35])
    wire mco_2_adj_610;   // mult_32s_2s.v(33[10:15])
    wire mult_32s_2s_0_mult_0_3_n1;   // mult_32s_2s.v(34[10:35])
    wire mult_32s_2s_0_mult_0_3_n0;   // mult_32s_2s.v(35[10:35])
    wire mco_3_adj_611;   // mult_32s_2s.v(38[10:15])
    wire mult_32s_2s_0_mult_0_4_n1;   // mult_32s_2s.v(39[10:35])
    wire mult_32s_2s_0_mult_0_4_n0;   // mult_32s_2s.v(40[10:35])
    wire mco_4_adj_612;   // mult_32s_2s.v(43[10:15])
    wire mult_32s_2s_0_mult_0_5_n1;   // mult_32s_2s.v(44[10:35])
    wire mult_32s_2s_0_mult_0_5_n0;   // mult_32s_2s.v(45[10:35])
    wire n73801 /* synthesis nomerge= */ ;
    
    wire n73840;
    wire [7:0]n1148;
    
    wire n23661, n63116, n63112, n63070, n63107, n63113, n63120, 
        n66804, n63130, n22437, n63114, n63150, n22106, n62900, 
        n22310, n41520, n62964, n25571, n73831, n39, n66628, n23655, 
        n23653, n63109, n23979, n23639;
    wire [27:0]n451_adj_700;
    wire [27:0]n480_adj_701;
    
    wire n63102;
    wire [7:0]n984;
    
    wire n63139, n63103;
    wire [27:0]n5;
    wire [27:0]n37_adj_763;
    
    wire n63111, n73809;
    wire [3:0]n3942;
    
    wire n3961, n15113;
    wire [63:0]n2022;
    wire [3:0]n1670;
    
    wire n73837;
    wire [7:0]n3980;
    
    wire n1682, n42934, n66796, n42939, n63156, n63068, n63104, 
        n63069, n63105, n63106, n63122, n63115, n27939, n73830, 
        n4599, n4617, n63147, n28181, n19214, n62966, n62961, 
        n66524, n66522, n24013, n63131, n23942, n23939, n73825, 
        n63128, n70867, n70866, n70855, n70835, n70834, n70833, 
        n62958, n70822, n66798, n70820, n70816, n35407, n73827, 
        n70788, n70778, n70771, n70744, n70740, n45598, n70727, 
        n73838, n63477, n66786, n70716, n73833, n73818, n67025, 
        n70693, n61382, n67007, n70692, n67005, n70691, n66961, 
        n66957, n66955;
    
    VHI i2 (.Z(inputNumber[2]));
    OSCH OSC0 (.STDBY(inputNumber[31]), .OSC(clock)) /* synthesis syn_instantiated=1 */ ;
    defparam OSC0.NOM_FREQ = "38.00";
    IB IBgsr (.I(GSRn), .O(GSRnX)) /* synthesis syn_black_box=true, syn_instantiated=1 */ ;
    GSR GSR_INST (.GSR(GSRnX)) /* synthesis syn_black_box=true, syn_noprune=true, syn_instantiated=1 */ ;
    BB BBspi_mosi (.I(spi_mosi_o), .T(spi_mosi_oe), .B(MOSI), .O(spi_mosi_i)) /* synthesis syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/spi.vhd(48[8:27])
    FADD2B mult_2u_2u_0_cin_lr_add_0 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_2u_2u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_3u_2u_0_cin_lr_add_0 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_3u_2u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_2u_3u_0_cin_lr_add_0 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_2u_3u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t7 (.A(A_int_adj_724[0]), .B(B_int_adj_725[8]), .Z(mult_24u_24u_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;
    FD1S1A dlatchrs_7_i2 (.D(writeout[1]), .CK(output_new), .Q(write_data[1]));
    defparam dlatchrs_7_i2.GSR = "DISABLED";
    FD1S1A dlatchrs_7_i3 (.D(writeout[2]), .CK(output_new), .Q(write_data[2]));
    defparam dlatchrs_7_i3.GSR = "DISABLED";
    FD1S1A dlatchrs_7_i4 (.D(writeout[3]), .CK(output_new), .Q(write_data[3]));
    defparam dlatchrs_7_i4.GSR = "DISABLED";
    FD1S1A dlatchrs_7_i5 (.D(writeout[4]), .CK(output_new), .Q(write_data[4]));
    defparam dlatchrs_7_i5.GSR = "DISABLED";
    FD1S1A dlatchrs_7_i6 (.D(writeout[5]), .CK(output_new), .Q(write_data[5]));
    defparam dlatchrs_7_i6.GSR = "DISABLED";
    FD1S1A dlatchrs_7_i7 (.D(writeout[6]), .CK(output_new), .Q(write_data[6]));
    defparam dlatchrs_7_i7.GSR = "DISABLED";
    FD1S1A dlatchrs_7_i8 (.D(writeout[7]), .CK(output_new), .Q(write_data[7]));
    defparam dlatchrs_7_i8.GSR = "DISABLED";
    BB BBspi_miso (.I(spi_miso_o), .T(spi_miso_oe), .B(MISO), .O(spi_miso_i)) /* synthesis syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/spi.vhd(48[8:27])
    BB BBspi_clk (.I(spi_clk_o), .T(spi_clk_oe), .B(SCLK), .O(spi_clk_i)) /* synthesis syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/spi.vhd(48[8:27])
    LUT4 m0_lut (.Z(n73801)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    LUT4 i53883_2_lut (.A(prod[35]), .B(prod[40]), .Z(n66786)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53883_2_lut.init = 16'heeee;
    LUT4 i53901_2_lut (.A(prod[32]), .B(prod[43]), .Z(n66804)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53901_2_lut.init = 16'heeee;
    LUT4 i54053_4_lut (.A(prod[46]), .B(prod[44]), .C(prod[33]), .D(prod[45]), 
         .Z(n66961)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54053_4_lut.init = 16'hfffe;
    LUT4 i53893_2_lut (.A(prod[22]), .B(prod[29]), .Z(n66796)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53893_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_801_4_lut (.A(B_int[7]), .B(A_int[7]), .C(diffExpAB[8]), 
         .D(diffExp[4]), .Z(n70771)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_801_4_lut.init = 16'hffca;
    LUT4 i54049_4_lut (.A(prod[42]), .B(prod[28]), .C(prod[41]), .D(prod[34]), 
         .Z(n66957)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54049_4_lut.init = 16'hfffe;
    LUT4 i53895_2_lut (.A(prod[24]), .B(prod[25]), .Z(n66798)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53895_2_lut.init = 16'heeee;
    LUT4 i54096_4_lut (.A(prod[27]), .B(n66961), .C(n66804), .D(prod[36]), 
         .Z(n67005)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54096_4_lut.init = 16'hfffe;
    LUT4 i24129_3_lut_rep_850 (.A(B_int[7]), .B(A_int[7]), .C(diffExpAB[8]), 
         .Z(n70820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24129_3_lut_rep_850.init = 16'hcaca;
    LUT4 i54098_4_lut (.A(n66786), .B(prod[38]), .C(prod[30]), .D(prod[39]), 
         .Z(n67007)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54098_4_lut.init = 16'hfffe;
    LUT4 i54114_4_lut (.A(n67005), .B(n66798), .C(n66957), .D(n66796), 
         .Z(n67025)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54114_4_lut.init = 16'hfffe;
    LUT4 i54047_4_lut (.A(prod[26]), .B(prod[37]), .C(prod[23]), .D(prod[31]), 
         .Z(n66955)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54047_4_lut.init = 16'hfffe;
    LUT4 i53916_4_lut (.A(n22437), .B(n25571), .C(n41520), .D(n22310), 
         .Z(n42934)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i53916_4_lut.init = 16'hfcdc;
    ND2 ND2_t31 (.A(i[1]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_0_n1)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_3u_2u_0_mult_0_1 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
          .A2(inputNumber[31]), .A3(inputNumber[31]), .B0(n70867), .B1(inputNumber[31]), 
          .B2(n70867), .B3(inputNumber[31]), .CI(mco_adj_572), .P0(n2889[3]), 
          .P1(n2889[4])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_3u_2u_0_mult_0_0 (.A0(inputNumber[2]), .A1(n14049[1]), .A2(n14049[1]), 
          .A3(inputNumber[31]), .B0(n70867), .B1(inputNumber[31]), .B2(n70867), 
          .B3(inputNumber[31]), .CI(mult_3u_2u_0_cin_lr_0), .CO(mco_adj_572), 
          .P0(n2889[1]), .P1(n2889[2])) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t0 (.A(inputNumber[2]), .B(inputNumber[31]), .Z(n2889[0])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_2u_2u_0_mult_0_0 (.A0(inputNumber[31]), .A1(n70867), .A2(n70867), 
          .A3(inputNumber[31]), .B0(n14049[1]), .B1(inputNumber[31]), 
          .B2(n14049[1]), .B3(inputNumber[31]), .CI(mult_2u_2u_0_cin_lr_0), 
          .CO(mfco_adj_573), .P0(n236[1]), .P1(n236[2])) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_2u_2u_0_Cadd_0_1 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_adj_573), 
           .S0(n236[3])) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t0_adj_983 (.A(inputNumber[31]), .B(inputNumber[31]), .Z(n236[0])) /* synthesis syn_instantiated=1 */ ;
    LUT4 mux_3895_i3_3_lut_rep_770_4_lut_4_lut (.A(diffExp[4]), .B(n70820), 
         .C(n70835), .D(n70833), .Z(n70740)) /* synthesis lut_function=(A (C+(D))+!A (B (C))) */ ;
    defparam mux_3895_i3_3_lut_rep_770_4_lut_4_lut.init = 16'heae0;
    LUT4 mux_3895_i11_4_lut_4_lut (.A(diffExp[4]), .B(n70820), .C(n70835), 
         .D(n70833), .Z(n37_adj_763[10])) /* synthesis lut_function=(!(A (C)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam mux_3895_i11_4_lut_4_lut.init = 16'h5e0e;
    AND2 AND2_t0_adj_984 (.A(inputNumber[2]), .B(inputNumber[31]), .Z(n3044[0])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_2u_3u_0_mult_0_0 (.A0(inputNumber[2]), .A1(n14053[1]), .A2(n14053[1]), 
          .A3(inputNumber[31]), .B0(n70867), .B1(inputNumber[31]), .B2(n70867), 
          .B3(inputNumber[31]), .CI(mult_2u_3u_0_cin_lr_0), .CO(mco_adj_571), 
          .P0(n3044[1]), .P1(n3044[2])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_2u_3u_0_mult_0_1 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
          .A2(inputNumber[31]), .A3(inputNumber[31]), .B0(n70867), .B1(inputNumber[31]), 
          .B2(n70867), .B3(inputNumber[31]), .CI(mco_adj_571), .P0(n3044[3]), 
          .P1(n3044[4])) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t8 (.A(A_int_adj_724[0]), .B(B_int_adj_725[6]), .Z(mult_24u_24u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t9 (.A(A_int_adj_724[0]), .B(B_int_adj_725[4]), .Z(mult_24u_24u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t10 (.A(A_int_adj_724[0]), .B(B_int_adj_725[2]), .Z(mult_24u_24u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_0_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco), .S0(mult_24u_24u_0_pp_0_25)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_2 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_2_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_1), .S0(mult_24u_24u_0_pp_1_27)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_4 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_4_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_2), .S0(mult_24u_24u_0_pp_2_29)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_6 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_6_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_3), .S0(mult_24u_24u_0_pp_3_31)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_8 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_8_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_4), .S0(mult_24u_24u_0_pp_4_33)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_10 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_10_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_5), .S0(mult_24u_24u_0_pp_5_35)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_12_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_6), .S0(mult_24u_24u_0_pp_6_37)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_14_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_7), .S0(mult_24u_24u_0_pp_7_39)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_16 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_16_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_8), .S0(mult_24u_24u_0_pp_8_41)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_18 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_18_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_9), .S0(mult_24u_24u_0_pp_9_43)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_20 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_20_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_10), .S0(mult_24u_24u_0_pp_10_45)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_22 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_Cadd_22_12 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(mfco_11), .S0(mult_24u_24u_0_pp_11_47)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_0_1 (.A0(inputNumber[31]), .A1(mult_24u_24u_0_pp_0_2), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_1_2), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_0_1)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_2 (.A0(mult_24u_24u_0_pp_0_3), .A1(mult_24u_24u_0_pp_0_4), 
           .B0(mult_24u_24u_0_pp_1_3), .B1(mult_24u_24u_0_pp_1_4), .CI(co_mult_24u_24u_0_0_1), 
           .COUT(co_mult_24u_24u_0_0_2), .S1(s_mult_24u_24u_0_0_4)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_3 (.A0(mult_24u_24u_0_pp_0_5), .A1(mult_24u_24u_0_pp_0_6), 
           .B0(mult_24u_24u_0_pp_1_5), .B1(mult_24u_24u_0_pp_1_6), .CI(co_mult_24u_24u_0_0_2), 
           .COUT(co_mult_24u_24u_0_0_3), .S0(s_mult_24u_24u_0_0_5), .S1(s_mult_24u_24u_0_0_6)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_4 (.A0(mult_24u_24u_0_pp_0_7), .A1(mult_24u_24u_0_pp_0_8), 
           .B0(mult_24u_24u_0_pp_1_7), .B1(mult_24u_24u_0_pp_1_8), .CI(co_mult_24u_24u_0_0_3), 
           .COUT(co_mult_24u_24u_0_0_4), .S0(s_mult_24u_24u_0_0_7), .S1(s_mult_24u_24u_0_0_8)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_5 (.A0(mult_24u_24u_0_pp_0_9), .A1(mult_24u_24u_0_pp_0_10), 
           .B0(mult_24u_24u_0_pp_1_9), .B1(mult_24u_24u_0_pp_1_10), .CI(co_mult_24u_24u_0_0_4), 
           .COUT(co_mult_24u_24u_0_0_5), .S0(s_mult_24u_24u_0_0_9), .S1(s_mult_24u_24u_0_0_10)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_6 (.A0(mult_24u_24u_0_pp_0_11), .A1(mult_24u_24u_0_pp_0_12), 
           .B0(mult_24u_24u_0_pp_1_11), .B1(mult_24u_24u_0_pp_1_12), .CI(co_mult_24u_24u_0_0_5), 
           .COUT(co_mult_24u_24u_0_0_6), .S0(s_mult_24u_24u_0_0_11), .S1(s_mult_24u_24u_0_0_12)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_7 (.A0(mult_24u_24u_0_pp_0_13), .A1(mult_24u_24u_0_pp_0_14), 
           .B0(mult_24u_24u_0_pp_1_13), .B1(mult_24u_24u_0_pp_1_14), .CI(co_mult_24u_24u_0_0_6), 
           .COUT(co_mult_24u_24u_0_0_7), .S0(s_mult_24u_24u_0_0_13), .S1(s_mult_24u_24u_0_0_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_8 (.A0(mult_24u_24u_0_pp_0_15), .A1(mult_24u_24u_0_pp_0_16), 
           .B0(mult_24u_24u_0_pp_1_15), .B1(mult_24u_24u_0_pp_1_16), .CI(co_mult_24u_24u_0_0_7), 
           .COUT(co_mult_24u_24u_0_0_8), .S0(s_mult_24u_24u_0_0_15), .S1(s_mult_24u_24u_0_0_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_9 (.A0(mult_24u_24u_0_pp_0_17), .A1(mult_24u_24u_0_pp_0_18), 
           .B0(mult_24u_24u_0_pp_1_17), .B1(mult_24u_24u_0_pp_1_18), .CI(co_mult_24u_24u_0_0_8), 
           .COUT(co_mult_24u_24u_0_0_9), .S0(s_mult_24u_24u_0_0_17), .S1(s_mult_24u_24u_0_0_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_10 (.A0(mult_24u_24u_0_pp_0_19), .A1(mult_24u_24u_0_pp_0_20), 
           .B0(mult_24u_24u_0_pp_1_19), .B1(mult_24u_24u_0_pp_1_20), .CI(co_mult_24u_24u_0_0_9), 
           .COUT(co_mult_24u_24u_0_0_10), .S0(s_mult_24u_24u_0_0_19), .S1(s_mult_24u_24u_0_0_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_11 (.A0(mult_24u_24u_0_pp_0_21), .A1(mult_24u_24u_0_pp_0_22), 
           .B0(mult_24u_24u_0_pp_1_21), .B1(mult_24u_24u_0_pp_1_22), .CI(co_mult_24u_24u_0_0_10), 
           .COUT(co_mult_24u_24u_0_0_11), .S0(s_mult_24u_24u_0_0_21), .S1(s_mult_24u_24u_0_0_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_12 (.A0(mult_24u_24u_0_pp_0_23), .A1(mult_24u_24u_0_pp_0_24), 
           .B0(mult_24u_24u_0_pp_1_23), .B1(mult_24u_24u_0_pp_1_24), .CI(co_mult_24u_24u_0_0_11), 
           .COUT(co_mult_24u_24u_0_0_12), .S0(s_mult_24u_24u_0_0_23), .S1(s_mult_24u_24u_0_0_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_13 (.A0(mult_24u_24u_0_pp_0_25), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_1_25), .B1(mult_24u_24u_0_pp_1_26), .CI(co_mult_24u_24u_0_0_12), 
           .COUT(co_mult_24u_24u_0_0_13), .S0(s_mult_24u_24u_0_0_25), .S1(s_mult_24u_24u_0_0_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_0_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_1_27), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_0_13), 
           .COUT(co_mult_24u_24u_0_0_14), .S0(s_mult_24u_24u_0_0_27), .S1(s_mult_24u_24u_0_0_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_0_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_0_14), 
           .S0(s_mult_24u_24u_0_0_29)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_1_1 (.A0(inputNumber[31]), .A1(mult_24u_24u_0_pp_2_6), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_3_6), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_1_1), .S1(s_mult_24u_24u_0_1_6)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_2 (.A0(mult_24u_24u_0_pp_2_7), .A1(mult_24u_24u_0_pp_2_8), 
           .B0(mult_24u_24u_0_pp_3_7), .B1(mult_24u_24u_0_pp_3_8), .CI(co_mult_24u_24u_0_1_1), 
           .COUT(co_mult_24u_24u_0_1_2), .S0(s_mult_24u_24u_0_1_7), .S1(s_mult_24u_24u_0_1_8)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_3 (.A0(mult_24u_24u_0_pp_2_9), .A1(mult_24u_24u_0_pp_2_10), 
           .B0(mult_24u_24u_0_pp_3_9), .B1(mult_24u_24u_0_pp_3_10), .CI(co_mult_24u_24u_0_1_2), 
           .COUT(co_mult_24u_24u_0_1_3), .S0(s_mult_24u_24u_0_1_9), .S1(s_mult_24u_24u_0_1_10)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_4 (.A0(mult_24u_24u_0_pp_2_11), .A1(mult_24u_24u_0_pp_2_12), 
           .B0(mult_24u_24u_0_pp_3_11), .B1(mult_24u_24u_0_pp_3_12), .CI(co_mult_24u_24u_0_1_3), 
           .COUT(co_mult_24u_24u_0_1_4), .S0(s_mult_24u_24u_0_1_11), .S1(s_mult_24u_24u_0_1_12)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_5 (.A0(mult_24u_24u_0_pp_2_13), .A1(mult_24u_24u_0_pp_2_14), 
           .B0(mult_24u_24u_0_pp_3_13), .B1(mult_24u_24u_0_pp_3_14), .CI(co_mult_24u_24u_0_1_4), 
           .COUT(co_mult_24u_24u_0_1_5), .S0(s_mult_24u_24u_0_1_13), .S1(s_mult_24u_24u_0_1_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_6 (.A0(mult_24u_24u_0_pp_2_15), .A1(mult_24u_24u_0_pp_2_16), 
           .B0(mult_24u_24u_0_pp_3_15), .B1(mult_24u_24u_0_pp_3_16), .CI(co_mult_24u_24u_0_1_5), 
           .COUT(co_mult_24u_24u_0_1_6), .S0(s_mult_24u_24u_0_1_15), .S1(s_mult_24u_24u_0_1_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_7 (.A0(mult_24u_24u_0_pp_2_17), .A1(mult_24u_24u_0_pp_2_18), 
           .B0(mult_24u_24u_0_pp_3_17), .B1(mult_24u_24u_0_pp_3_18), .CI(co_mult_24u_24u_0_1_6), 
           .COUT(co_mult_24u_24u_0_1_7), .S0(s_mult_24u_24u_0_1_17), .S1(s_mult_24u_24u_0_1_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_8 (.A0(mult_24u_24u_0_pp_2_19), .A1(mult_24u_24u_0_pp_2_20), 
           .B0(mult_24u_24u_0_pp_3_19), .B1(mult_24u_24u_0_pp_3_20), .CI(co_mult_24u_24u_0_1_7), 
           .COUT(co_mult_24u_24u_0_1_8), .S0(s_mult_24u_24u_0_1_19), .S1(s_mult_24u_24u_0_1_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_9 (.A0(mult_24u_24u_0_pp_2_21), .A1(mult_24u_24u_0_pp_2_22), 
           .B0(mult_24u_24u_0_pp_3_21), .B1(mult_24u_24u_0_pp_3_22), .CI(co_mult_24u_24u_0_1_8), 
           .COUT(co_mult_24u_24u_0_1_9), .S0(s_mult_24u_24u_0_1_21), .S1(s_mult_24u_24u_0_1_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_10 (.A0(mult_24u_24u_0_pp_2_23), .A1(mult_24u_24u_0_pp_2_24), 
           .B0(mult_24u_24u_0_pp_3_23), .B1(mult_24u_24u_0_pp_3_24), .CI(co_mult_24u_24u_0_1_9), 
           .COUT(co_mult_24u_24u_0_1_10), .S0(s_mult_24u_24u_0_1_23), .S1(s_mult_24u_24u_0_1_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_11 (.A0(mult_24u_24u_0_pp_2_25), .A1(mult_24u_24u_0_pp_2_26), 
           .B0(mult_24u_24u_0_pp_3_25), .B1(mult_24u_24u_0_pp_3_26), .CI(co_mult_24u_24u_0_1_10), 
           .COUT(co_mult_24u_24u_0_1_11), .S0(s_mult_24u_24u_0_1_25), .S1(s_mult_24u_24u_0_1_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_12 (.A0(mult_24u_24u_0_pp_2_27), .A1(mult_24u_24u_0_pp_2_28), 
           .B0(mult_24u_24u_0_pp_3_27), .B1(mult_24u_24u_0_pp_3_28), .CI(co_mult_24u_24u_0_1_11), 
           .COUT(co_mult_24u_24u_0_1_12), .S0(s_mult_24u_24u_0_1_27), .S1(s_mult_24u_24u_0_1_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_13 (.A0(mult_24u_24u_0_pp_2_29), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_3_29), .B1(mult_24u_24u_0_pp_3_30), .CI(co_mult_24u_24u_0_1_12), 
           .COUT(co_mult_24u_24u_0_1_13), .S0(s_mult_24u_24u_0_1_29), .S1(s_mult_24u_24u_0_1_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_1_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_3_31), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_1_13), 
           .COUT(co_mult_24u_24u_0_1_14), .S0(s_mult_24u_24u_0_1_31), .S1(s_mult_24u_24u_0_1_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_1_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_1_14), 
           .S0(s_mult_24u_24u_0_1_33)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_2_1 (.A0(inputNumber[31]), .A1(mult_24u_24u_0_pp_4_10), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_5_10), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_2_1), .S1(s_mult_24u_24u_0_2_10)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_2 (.A0(mult_24u_24u_0_pp_4_11), .A1(mult_24u_24u_0_pp_4_12), 
           .B0(mult_24u_24u_0_pp_5_11), .B1(mult_24u_24u_0_pp_5_12), .CI(co_mult_24u_24u_0_2_1), 
           .COUT(co_mult_24u_24u_0_2_2), .S0(s_mult_24u_24u_0_2_11), .S1(s_mult_24u_24u_0_2_12)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_3 (.A0(mult_24u_24u_0_pp_4_13), .A1(mult_24u_24u_0_pp_4_14), 
           .B0(mult_24u_24u_0_pp_5_13), .B1(mult_24u_24u_0_pp_5_14), .CI(co_mult_24u_24u_0_2_2), 
           .COUT(co_mult_24u_24u_0_2_3), .S0(s_mult_24u_24u_0_2_13), .S1(s_mult_24u_24u_0_2_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_4 (.A0(mult_24u_24u_0_pp_4_15), .A1(mult_24u_24u_0_pp_4_16), 
           .B0(mult_24u_24u_0_pp_5_15), .B1(mult_24u_24u_0_pp_5_16), .CI(co_mult_24u_24u_0_2_3), 
           .COUT(co_mult_24u_24u_0_2_4), .S0(s_mult_24u_24u_0_2_15), .S1(s_mult_24u_24u_0_2_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_5 (.A0(mult_24u_24u_0_pp_4_17), .A1(mult_24u_24u_0_pp_4_18), 
           .B0(mult_24u_24u_0_pp_5_17), .B1(mult_24u_24u_0_pp_5_18), .CI(co_mult_24u_24u_0_2_4), 
           .COUT(co_mult_24u_24u_0_2_5), .S0(s_mult_24u_24u_0_2_17), .S1(s_mult_24u_24u_0_2_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_6 (.A0(mult_24u_24u_0_pp_4_19), .A1(mult_24u_24u_0_pp_4_20), 
           .B0(mult_24u_24u_0_pp_5_19), .B1(mult_24u_24u_0_pp_5_20), .CI(co_mult_24u_24u_0_2_5), 
           .COUT(co_mult_24u_24u_0_2_6), .S0(s_mult_24u_24u_0_2_19), .S1(s_mult_24u_24u_0_2_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_7 (.A0(mult_24u_24u_0_pp_4_21), .A1(mult_24u_24u_0_pp_4_22), 
           .B0(mult_24u_24u_0_pp_5_21), .B1(mult_24u_24u_0_pp_5_22), .CI(co_mult_24u_24u_0_2_6), 
           .COUT(co_mult_24u_24u_0_2_7), .S0(s_mult_24u_24u_0_2_21), .S1(s_mult_24u_24u_0_2_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_8 (.A0(mult_24u_24u_0_pp_4_23), .A1(mult_24u_24u_0_pp_4_24), 
           .B0(mult_24u_24u_0_pp_5_23), .B1(mult_24u_24u_0_pp_5_24), .CI(co_mult_24u_24u_0_2_7), 
           .COUT(co_mult_24u_24u_0_2_8), .S0(s_mult_24u_24u_0_2_23), .S1(s_mult_24u_24u_0_2_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_9 (.A0(mult_24u_24u_0_pp_4_25), .A1(mult_24u_24u_0_pp_4_26), 
           .B0(mult_24u_24u_0_pp_5_25), .B1(mult_24u_24u_0_pp_5_26), .CI(co_mult_24u_24u_0_2_8), 
           .COUT(co_mult_24u_24u_0_2_9), .S0(s_mult_24u_24u_0_2_25), .S1(s_mult_24u_24u_0_2_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_10 (.A0(mult_24u_24u_0_pp_4_27), .A1(mult_24u_24u_0_pp_4_28), 
           .B0(mult_24u_24u_0_pp_5_27), .B1(mult_24u_24u_0_pp_5_28), .CI(co_mult_24u_24u_0_2_9), 
           .COUT(co_mult_24u_24u_0_2_10), .S0(s_mult_24u_24u_0_2_27), .S1(s_mult_24u_24u_0_2_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_11 (.A0(mult_24u_24u_0_pp_4_29), .A1(mult_24u_24u_0_pp_4_30), 
           .B0(mult_24u_24u_0_pp_5_29), .B1(mult_24u_24u_0_pp_5_30), .CI(co_mult_24u_24u_0_2_10), 
           .COUT(co_mult_24u_24u_0_2_11), .S0(s_mult_24u_24u_0_2_29), .S1(s_mult_24u_24u_0_2_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_12 (.A0(mult_24u_24u_0_pp_4_31), .A1(mult_24u_24u_0_pp_4_32), 
           .B0(mult_24u_24u_0_pp_5_31), .B1(mult_24u_24u_0_pp_5_32), .CI(co_mult_24u_24u_0_2_11), 
           .COUT(co_mult_24u_24u_0_2_12), .S0(s_mult_24u_24u_0_2_31), .S1(s_mult_24u_24u_0_2_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_13 (.A0(mult_24u_24u_0_pp_4_33), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_5_33), .B1(mult_24u_24u_0_pp_5_34), .CI(co_mult_24u_24u_0_2_12), 
           .COUT(co_mult_24u_24u_0_2_13), .S0(s_mult_24u_24u_0_2_33), .S1(s_mult_24u_24u_0_2_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_2_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_5_35), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_2_13), 
           .COUT(co_mult_24u_24u_0_2_14), .S0(s_mult_24u_24u_0_2_35), .S1(s_mult_24u_24u_0_2_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_2_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_2_14), 
           .S0(s_mult_24u_24u_0_2_37)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_3_1 (.A0(inputNumber[31]), .A1(mult_24u_24u_0_pp_6_14), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_7_14), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_3_1), .S1(s_mult_24u_24u_0_3_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_2 (.A0(mult_24u_24u_0_pp_6_15), .A1(mult_24u_24u_0_pp_6_16), 
           .B0(mult_24u_24u_0_pp_7_15), .B1(mult_24u_24u_0_pp_7_16), .CI(co_mult_24u_24u_0_3_1), 
           .COUT(co_mult_24u_24u_0_3_2), .S0(s_mult_24u_24u_0_3_15), .S1(s_mult_24u_24u_0_3_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_3 (.A0(mult_24u_24u_0_pp_6_17), .A1(mult_24u_24u_0_pp_6_18), 
           .B0(mult_24u_24u_0_pp_7_17), .B1(mult_24u_24u_0_pp_7_18), .CI(co_mult_24u_24u_0_3_2), 
           .COUT(co_mult_24u_24u_0_3_3), .S0(s_mult_24u_24u_0_3_17), .S1(s_mult_24u_24u_0_3_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_4 (.A0(mult_24u_24u_0_pp_6_19), .A1(mult_24u_24u_0_pp_6_20), 
           .B0(mult_24u_24u_0_pp_7_19), .B1(mult_24u_24u_0_pp_7_20), .CI(co_mult_24u_24u_0_3_3), 
           .COUT(co_mult_24u_24u_0_3_4), .S0(s_mult_24u_24u_0_3_19), .S1(s_mult_24u_24u_0_3_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_5 (.A0(mult_24u_24u_0_pp_6_21), .A1(mult_24u_24u_0_pp_6_22), 
           .B0(mult_24u_24u_0_pp_7_21), .B1(mult_24u_24u_0_pp_7_22), .CI(co_mult_24u_24u_0_3_4), 
           .COUT(co_mult_24u_24u_0_3_5), .S0(s_mult_24u_24u_0_3_21), .S1(s_mult_24u_24u_0_3_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_6 (.A0(mult_24u_24u_0_pp_6_23), .A1(mult_24u_24u_0_pp_6_24), 
           .B0(mult_24u_24u_0_pp_7_23), .B1(mult_24u_24u_0_pp_7_24), .CI(co_mult_24u_24u_0_3_5), 
           .COUT(co_mult_24u_24u_0_3_6), .S0(s_mult_24u_24u_0_3_23), .S1(s_mult_24u_24u_0_3_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_7 (.A0(mult_24u_24u_0_pp_6_25), .A1(mult_24u_24u_0_pp_6_26), 
           .B0(mult_24u_24u_0_pp_7_25), .B1(mult_24u_24u_0_pp_7_26), .CI(co_mult_24u_24u_0_3_6), 
           .COUT(co_mult_24u_24u_0_3_7), .S0(s_mult_24u_24u_0_3_25), .S1(s_mult_24u_24u_0_3_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_8 (.A0(mult_24u_24u_0_pp_6_27), .A1(mult_24u_24u_0_pp_6_28), 
           .B0(mult_24u_24u_0_pp_7_27), .B1(mult_24u_24u_0_pp_7_28), .CI(co_mult_24u_24u_0_3_7), 
           .COUT(co_mult_24u_24u_0_3_8), .S0(s_mult_24u_24u_0_3_27), .S1(s_mult_24u_24u_0_3_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_9 (.A0(mult_24u_24u_0_pp_6_29), .A1(mult_24u_24u_0_pp_6_30), 
           .B0(mult_24u_24u_0_pp_7_29), .B1(mult_24u_24u_0_pp_7_30), .CI(co_mult_24u_24u_0_3_8), 
           .COUT(co_mult_24u_24u_0_3_9), .S0(s_mult_24u_24u_0_3_29), .S1(s_mult_24u_24u_0_3_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_10 (.A0(mult_24u_24u_0_pp_6_31), .A1(mult_24u_24u_0_pp_6_32), 
           .B0(mult_24u_24u_0_pp_7_31), .B1(mult_24u_24u_0_pp_7_32), .CI(co_mult_24u_24u_0_3_9), 
           .COUT(co_mult_24u_24u_0_3_10), .S0(s_mult_24u_24u_0_3_31), .S1(s_mult_24u_24u_0_3_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_11 (.A0(mult_24u_24u_0_pp_6_33), .A1(mult_24u_24u_0_pp_6_34), 
           .B0(mult_24u_24u_0_pp_7_33), .B1(mult_24u_24u_0_pp_7_34), .CI(co_mult_24u_24u_0_3_10), 
           .COUT(co_mult_24u_24u_0_3_11), .S0(s_mult_24u_24u_0_3_33), .S1(s_mult_24u_24u_0_3_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_12 (.A0(mult_24u_24u_0_pp_6_35), .A1(mult_24u_24u_0_pp_6_36), 
           .B0(mult_24u_24u_0_pp_7_35), .B1(mult_24u_24u_0_pp_7_36), .CI(co_mult_24u_24u_0_3_11), 
           .COUT(co_mult_24u_24u_0_3_12), .S0(s_mult_24u_24u_0_3_35), .S1(s_mult_24u_24u_0_3_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_13 (.A0(mult_24u_24u_0_pp_6_37), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_7_37), .B1(mult_24u_24u_0_pp_7_38), .CI(co_mult_24u_24u_0_3_12), 
           .COUT(co_mult_24u_24u_0_3_13), .S0(s_mult_24u_24u_0_3_37), .S1(s_mult_24u_24u_0_3_38)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_3_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_7_39), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_3_13), 
           .COUT(co_mult_24u_24u_0_3_14), .S0(s_mult_24u_24u_0_3_39), .S1(s_mult_24u_24u_0_3_40)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_3_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_3_14), 
           .S0(s_mult_24u_24u_0_3_41)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_4_1 (.A0(inputNumber[31]), .A1(mult_24u_24u_0_pp_8_18), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_9_18), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_4_1), .S1(s_mult_24u_24u_0_4_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_2 (.A0(mult_24u_24u_0_pp_8_19), .A1(mult_24u_24u_0_pp_8_20), 
           .B0(mult_24u_24u_0_pp_9_19), .B1(mult_24u_24u_0_pp_9_20), .CI(co_mult_24u_24u_0_4_1), 
           .COUT(co_mult_24u_24u_0_4_2), .S0(s_mult_24u_24u_0_4_19), .S1(s_mult_24u_24u_0_4_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_3 (.A0(mult_24u_24u_0_pp_8_21), .A1(mult_24u_24u_0_pp_8_22), 
           .B0(mult_24u_24u_0_pp_9_21), .B1(mult_24u_24u_0_pp_9_22), .CI(co_mult_24u_24u_0_4_2), 
           .COUT(co_mult_24u_24u_0_4_3), .S0(s_mult_24u_24u_0_4_21), .S1(s_mult_24u_24u_0_4_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_4 (.A0(mult_24u_24u_0_pp_8_23), .A1(mult_24u_24u_0_pp_8_24), 
           .B0(mult_24u_24u_0_pp_9_23), .B1(mult_24u_24u_0_pp_9_24), .CI(co_mult_24u_24u_0_4_3), 
           .COUT(co_mult_24u_24u_0_4_4), .S0(s_mult_24u_24u_0_4_23), .S1(s_mult_24u_24u_0_4_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_5 (.A0(mult_24u_24u_0_pp_8_25), .A1(mult_24u_24u_0_pp_8_26), 
           .B0(mult_24u_24u_0_pp_9_25), .B1(mult_24u_24u_0_pp_9_26), .CI(co_mult_24u_24u_0_4_4), 
           .COUT(co_mult_24u_24u_0_4_5), .S0(s_mult_24u_24u_0_4_25), .S1(s_mult_24u_24u_0_4_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_6 (.A0(mult_24u_24u_0_pp_8_27), .A1(mult_24u_24u_0_pp_8_28), 
           .B0(mult_24u_24u_0_pp_9_27), .B1(mult_24u_24u_0_pp_9_28), .CI(co_mult_24u_24u_0_4_5), 
           .COUT(co_mult_24u_24u_0_4_6), .S0(s_mult_24u_24u_0_4_27), .S1(s_mult_24u_24u_0_4_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_7 (.A0(mult_24u_24u_0_pp_8_29), .A1(mult_24u_24u_0_pp_8_30), 
           .B0(mult_24u_24u_0_pp_9_29), .B1(mult_24u_24u_0_pp_9_30), .CI(co_mult_24u_24u_0_4_6), 
           .COUT(co_mult_24u_24u_0_4_7), .S0(s_mult_24u_24u_0_4_29), .S1(s_mult_24u_24u_0_4_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_8 (.A0(mult_24u_24u_0_pp_8_31), .A1(mult_24u_24u_0_pp_8_32), 
           .B0(mult_24u_24u_0_pp_9_31), .B1(mult_24u_24u_0_pp_9_32), .CI(co_mult_24u_24u_0_4_7), 
           .COUT(co_mult_24u_24u_0_4_8), .S0(s_mult_24u_24u_0_4_31), .S1(s_mult_24u_24u_0_4_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_9 (.A0(mult_24u_24u_0_pp_8_33), .A1(mult_24u_24u_0_pp_8_34), 
           .B0(mult_24u_24u_0_pp_9_33), .B1(mult_24u_24u_0_pp_9_34), .CI(co_mult_24u_24u_0_4_8), 
           .COUT(co_mult_24u_24u_0_4_9), .S0(s_mult_24u_24u_0_4_33), .S1(s_mult_24u_24u_0_4_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_10 (.A0(mult_24u_24u_0_pp_8_35), .A1(mult_24u_24u_0_pp_8_36), 
           .B0(mult_24u_24u_0_pp_9_35), .B1(mult_24u_24u_0_pp_9_36), .CI(co_mult_24u_24u_0_4_9), 
           .COUT(co_mult_24u_24u_0_4_10), .S0(s_mult_24u_24u_0_4_35), .S1(s_mult_24u_24u_0_4_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_11 (.A0(mult_24u_24u_0_pp_8_37), .A1(mult_24u_24u_0_pp_8_38), 
           .B0(mult_24u_24u_0_pp_9_37), .B1(mult_24u_24u_0_pp_9_38), .CI(co_mult_24u_24u_0_4_10), 
           .COUT(co_mult_24u_24u_0_4_11), .S0(s_mult_24u_24u_0_4_37), .S1(s_mult_24u_24u_0_4_38)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_12 (.A0(mult_24u_24u_0_pp_8_39), .A1(mult_24u_24u_0_pp_8_40), 
           .B0(mult_24u_24u_0_pp_9_39), .B1(mult_24u_24u_0_pp_9_40), .CI(co_mult_24u_24u_0_4_11), 
           .COUT(co_mult_24u_24u_0_4_12), .S0(s_mult_24u_24u_0_4_39), .S1(s_mult_24u_24u_0_4_40)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_13 (.A0(mult_24u_24u_0_pp_8_41), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_9_41), .B1(mult_24u_24u_0_pp_9_42), .CI(co_mult_24u_24u_0_4_12), 
           .COUT(co_mult_24u_24u_0_4_13), .S0(s_mult_24u_24u_0_4_41), .S1(s_mult_24u_24u_0_4_42)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_4_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_9_43), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_4_13), 
           .COUT(co_mult_24u_24u_0_4_14), .S0(s_mult_24u_24u_0_4_43), .S1(s_mult_24u_24u_0_4_44)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_4_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_4_14), 
           .S0(s_mult_24u_24u_0_4_45)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_5_1 (.A0(inputNumber[31]), .A1(mult_24u_24u_0_pp_10_22), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_11_22), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_5_1), .S1(s_mult_24u_24u_0_5_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_2 (.A0(mult_24u_24u_0_pp_10_23), .A1(mult_24u_24u_0_pp_10_24), 
           .B0(mult_24u_24u_0_pp_11_23), .B1(mult_24u_24u_0_pp_11_24), .CI(co_mult_24u_24u_0_5_1), 
           .COUT(co_mult_24u_24u_0_5_2), .S0(s_mult_24u_24u_0_5_23), .S1(s_mult_24u_24u_0_5_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_3 (.A0(mult_24u_24u_0_pp_10_25), .A1(mult_24u_24u_0_pp_10_26), 
           .B0(mult_24u_24u_0_pp_11_25), .B1(mult_24u_24u_0_pp_11_26), .CI(co_mult_24u_24u_0_5_2), 
           .COUT(co_mult_24u_24u_0_5_3), .S0(s_mult_24u_24u_0_5_25), .S1(s_mult_24u_24u_0_5_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_4 (.A0(mult_24u_24u_0_pp_10_27), .A1(mult_24u_24u_0_pp_10_28), 
           .B0(mult_24u_24u_0_pp_11_27), .B1(mult_24u_24u_0_pp_11_28), .CI(co_mult_24u_24u_0_5_3), 
           .COUT(co_mult_24u_24u_0_5_4), .S0(s_mult_24u_24u_0_5_27), .S1(s_mult_24u_24u_0_5_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_5 (.A0(mult_24u_24u_0_pp_10_29), .A1(mult_24u_24u_0_pp_10_30), 
           .B0(mult_24u_24u_0_pp_11_29), .B1(mult_24u_24u_0_pp_11_30), .CI(co_mult_24u_24u_0_5_4), 
           .COUT(co_mult_24u_24u_0_5_5), .S0(s_mult_24u_24u_0_5_29), .S1(s_mult_24u_24u_0_5_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_6 (.A0(mult_24u_24u_0_pp_10_31), .A1(mult_24u_24u_0_pp_10_32), 
           .B0(mult_24u_24u_0_pp_11_31), .B1(mult_24u_24u_0_pp_11_32), .CI(co_mult_24u_24u_0_5_5), 
           .COUT(co_mult_24u_24u_0_5_6), .S0(s_mult_24u_24u_0_5_31), .S1(s_mult_24u_24u_0_5_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_7 (.A0(mult_24u_24u_0_pp_10_33), .A1(mult_24u_24u_0_pp_10_34), 
           .B0(mult_24u_24u_0_pp_11_33), .B1(mult_24u_24u_0_pp_11_34), .CI(co_mult_24u_24u_0_5_6), 
           .COUT(co_mult_24u_24u_0_5_7), .S0(s_mult_24u_24u_0_5_33), .S1(s_mult_24u_24u_0_5_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_8 (.A0(mult_24u_24u_0_pp_10_35), .A1(mult_24u_24u_0_pp_10_36), 
           .B0(mult_24u_24u_0_pp_11_35), .B1(mult_24u_24u_0_pp_11_36), .CI(co_mult_24u_24u_0_5_7), 
           .COUT(co_mult_24u_24u_0_5_8), .S0(s_mult_24u_24u_0_5_35), .S1(s_mult_24u_24u_0_5_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_9 (.A0(mult_24u_24u_0_pp_10_37), .A1(mult_24u_24u_0_pp_10_38), 
           .B0(mult_24u_24u_0_pp_11_37), .B1(mult_24u_24u_0_pp_11_38), .CI(co_mult_24u_24u_0_5_8), 
           .COUT(co_mult_24u_24u_0_5_9), .S0(s_mult_24u_24u_0_5_37), .S1(s_mult_24u_24u_0_5_38)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_10 (.A0(mult_24u_24u_0_pp_10_39), .A1(mult_24u_24u_0_pp_10_40), 
           .B0(mult_24u_24u_0_pp_11_39), .B1(mult_24u_24u_0_pp_11_40), .CI(co_mult_24u_24u_0_5_9), 
           .COUT(co_mult_24u_24u_0_5_10), .S0(s_mult_24u_24u_0_5_39), .S1(s_mult_24u_24u_0_5_40)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_11 (.A0(mult_24u_24u_0_pp_10_41), .A1(mult_24u_24u_0_pp_10_42), 
           .B0(mult_24u_24u_0_pp_11_41), .B1(mult_24u_24u_0_pp_11_42), .CI(co_mult_24u_24u_0_5_10), 
           .COUT(co_mult_24u_24u_0_5_11), .S0(s_mult_24u_24u_0_5_41), .S1(s_mult_24u_24u_0_5_42)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_12 (.A0(mult_24u_24u_0_pp_10_43), .A1(mult_24u_24u_0_pp_10_44), 
           .B0(mult_24u_24u_0_pp_11_43), .B1(mult_24u_24u_0_pp_11_44), .CI(co_mult_24u_24u_0_5_11), 
           .COUT(co_mult_24u_24u_0_5_12), .S0(s_mult_24u_24u_0_5_43), .S1(s_mult_24u_24u_0_5_44)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_13 (.A0(mult_24u_24u_0_pp_10_45), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_11_45), .B1(mult_24u_24u_0_pp_11_46), .CI(co_mult_24u_24u_0_5_12), 
           .COUT(co_mult_24u_24u_0_5_13), .S0(s_mult_24u_24u_0_5_45), .S1(s_mult_24u_24u_0_5_46)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_5_14 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(mult_24u_24u_0_pp_11_47), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_5_13), 
           .S0(s_mult_24u_24u_0_5_47)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_6_1 (.A0(inputNumber[31]), .A1(s_mult_24u_24u_0_0_4), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_2_4), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_6_1)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_2 (.A0(s_mult_24u_24u_0_0_5), .A1(s_mult_24u_24u_0_0_6), 
           .B0(mult_24u_24u_0_pp_2_5), .B1(s_mult_24u_24u_0_1_6), .CI(co_mult_24u_24u_0_6_1), 
           .COUT(co_mult_24u_24u_0_6_2)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_3 (.A0(s_mult_24u_24u_0_0_7), .A1(s_mult_24u_24u_0_0_8), 
           .B0(s_mult_24u_24u_0_1_7), .B1(s_mult_24u_24u_0_1_8), .CI(co_mult_24u_24u_0_6_2), 
           .COUT(co_mult_24u_24u_0_6_3), .S1(s_mult_24u_24u_0_6_8)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_4 (.A0(s_mult_24u_24u_0_0_9), .A1(s_mult_24u_24u_0_0_10), 
           .B0(s_mult_24u_24u_0_1_9), .B1(s_mult_24u_24u_0_1_10), .CI(co_mult_24u_24u_0_6_3), 
           .COUT(co_mult_24u_24u_0_6_4), .S0(s_mult_24u_24u_0_6_9), .S1(s_mult_24u_24u_0_6_10)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_5 (.A0(s_mult_24u_24u_0_0_11), .A1(s_mult_24u_24u_0_0_12), 
           .B0(s_mult_24u_24u_0_1_11), .B1(s_mult_24u_24u_0_1_12), .CI(co_mult_24u_24u_0_6_4), 
           .COUT(co_mult_24u_24u_0_6_5), .S0(s_mult_24u_24u_0_6_11), .S1(s_mult_24u_24u_0_6_12)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_6 (.A0(s_mult_24u_24u_0_0_13), .A1(s_mult_24u_24u_0_0_14), 
           .B0(s_mult_24u_24u_0_1_13), .B1(s_mult_24u_24u_0_1_14), .CI(co_mult_24u_24u_0_6_5), 
           .COUT(co_mult_24u_24u_0_6_6), .S0(s_mult_24u_24u_0_6_13), .S1(s_mult_24u_24u_0_6_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_7 (.A0(s_mult_24u_24u_0_0_15), .A1(s_mult_24u_24u_0_0_16), 
           .B0(s_mult_24u_24u_0_1_15), .B1(s_mult_24u_24u_0_1_16), .CI(co_mult_24u_24u_0_6_6), 
           .COUT(co_mult_24u_24u_0_6_7), .S0(s_mult_24u_24u_0_6_15), .S1(s_mult_24u_24u_0_6_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_8 (.A0(s_mult_24u_24u_0_0_17), .A1(s_mult_24u_24u_0_0_18), 
           .B0(s_mult_24u_24u_0_1_17), .B1(s_mult_24u_24u_0_1_18), .CI(co_mult_24u_24u_0_6_7), 
           .COUT(co_mult_24u_24u_0_6_8), .S0(s_mult_24u_24u_0_6_17), .S1(s_mult_24u_24u_0_6_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_9 (.A0(s_mult_24u_24u_0_0_19), .A1(s_mult_24u_24u_0_0_20), 
           .B0(s_mult_24u_24u_0_1_19), .B1(s_mult_24u_24u_0_1_20), .CI(co_mult_24u_24u_0_6_8), 
           .COUT(co_mult_24u_24u_0_6_9), .S0(s_mult_24u_24u_0_6_19), .S1(s_mult_24u_24u_0_6_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_10 (.A0(s_mult_24u_24u_0_0_21), .A1(s_mult_24u_24u_0_0_22), 
           .B0(s_mult_24u_24u_0_1_21), .B1(s_mult_24u_24u_0_1_22), .CI(co_mult_24u_24u_0_6_9), 
           .COUT(co_mult_24u_24u_0_6_10), .S0(s_mult_24u_24u_0_6_21), .S1(s_mult_24u_24u_0_6_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_11 (.A0(s_mult_24u_24u_0_0_23), .A1(s_mult_24u_24u_0_0_24), 
           .B0(s_mult_24u_24u_0_1_23), .B1(s_mult_24u_24u_0_1_24), .CI(co_mult_24u_24u_0_6_10), 
           .COUT(co_mult_24u_24u_0_6_11), .S0(s_mult_24u_24u_0_6_23), .S1(s_mult_24u_24u_0_6_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_12 (.A0(s_mult_24u_24u_0_0_25), .A1(s_mult_24u_24u_0_0_26), 
           .B0(s_mult_24u_24u_0_1_25), .B1(s_mult_24u_24u_0_1_26), .CI(co_mult_24u_24u_0_6_11), 
           .COUT(co_mult_24u_24u_0_6_12), .S0(s_mult_24u_24u_0_6_25), .S1(s_mult_24u_24u_0_6_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_13 (.A0(s_mult_24u_24u_0_0_27), .A1(s_mult_24u_24u_0_0_28), 
           .B0(s_mult_24u_24u_0_1_27), .B1(s_mult_24u_24u_0_1_28), .CI(co_mult_24u_24u_0_6_12), 
           .COUT(co_mult_24u_24u_0_6_13), .S0(s_mult_24u_24u_0_6_27), .S1(s_mult_24u_24u_0_6_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_14 (.A0(s_mult_24u_24u_0_0_29), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_1_29), .B1(s_mult_24u_24u_0_1_30), .CI(co_mult_24u_24u_0_6_13), 
           .COUT(co_mult_24u_24u_0_6_14), .S0(s_mult_24u_24u_0_6_29), .S1(s_mult_24u_24u_0_6_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_1_31), .B1(s_mult_24u_24u_0_1_32), .CI(co_mult_24u_24u_0_6_14), 
           .COUT(co_mult_24u_24u_0_6_15), .S0(s_mult_24u_24u_0_6_31), .S1(s_mult_24u_24u_0_6_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_6_16 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_1_33), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_6_15), 
           .COUT(co_mult_24u_24u_0_6_16), .S0(s_mult_24u_24u_0_6_33), .S1(s_mult_24u_24u_0_6_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_6_17 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_6_16), 
           .S0(s_mult_24u_24u_0_6_35)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_7_1 (.A0(inputNumber[31]), .A1(s_mult_24u_24u_0_2_12), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_6_12), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_7_1), .S1(s_mult_24u_24u_0_7_12)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_2 (.A0(s_mult_24u_24u_0_2_13), .A1(s_mult_24u_24u_0_2_14), 
           .B0(mult_24u_24u_0_pp_6_13), .B1(s_mult_24u_24u_0_3_14), .CI(co_mult_24u_24u_0_7_1), 
           .COUT(co_mult_24u_24u_0_7_2), .S0(s_mult_24u_24u_0_7_13), .S1(s_mult_24u_24u_0_7_14)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_3 (.A0(s_mult_24u_24u_0_2_15), .A1(s_mult_24u_24u_0_2_16), 
           .B0(s_mult_24u_24u_0_3_15), .B1(s_mult_24u_24u_0_3_16), .CI(co_mult_24u_24u_0_7_2), 
           .COUT(co_mult_24u_24u_0_7_3), .S0(s_mult_24u_24u_0_7_15), .S1(s_mult_24u_24u_0_7_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_4 (.A0(s_mult_24u_24u_0_2_17), .A1(s_mult_24u_24u_0_2_18), 
           .B0(s_mult_24u_24u_0_3_17), .B1(s_mult_24u_24u_0_3_18), .CI(co_mult_24u_24u_0_7_3), 
           .COUT(co_mult_24u_24u_0_7_4), .S0(s_mult_24u_24u_0_7_17), .S1(s_mult_24u_24u_0_7_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_5 (.A0(s_mult_24u_24u_0_2_19), .A1(s_mult_24u_24u_0_2_20), 
           .B0(s_mult_24u_24u_0_3_19), .B1(s_mult_24u_24u_0_3_20), .CI(co_mult_24u_24u_0_7_4), 
           .COUT(co_mult_24u_24u_0_7_5), .S0(s_mult_24u_24u_0_7_19), .S1(s_mult_24u_24u_0_7_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_6 (.A0(s_mult_24u_24u_0_2_21), .A1(s_mult_24u_24u_0_2_22), 
           .B0(s_mult_24u_24u_0_3_21), .B1(s_mult_24u_24u_0_3_22), .CI(co_mult_24u_24u_0_7_5), 
           .COUT(co_mult_24u_24u_0_7_6), .S0(s_mult_24u_24u_0_7_21), .S1(s_mult_24u_24u_0_7_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_7 (.A0(s_mult_24u_24u_0_2_23), .A1(s_mult_24u_24u_0_2_24), 
           .B0(s_mult_24u_24u_0_3_23), .B1(s_mult_24u_24u_0_3_24), .CI(co_mult_24u_24u_0_7_6), 
           .COUT(co_mult_24u_24u_0_7_7), .S0(s_mult_24u_24u_0_7_23), .S1(s_mult_24u_24u_0_7_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_8 (.A0(s_mult_24u_24u_0_2_25), .A1(s_mult_24u_24u_0_2_26), 
           .B0(s_mult_24u_24u_0_3_25), .B1(s_mult_24u_24u_0_3_26), .CI(co_mult_24u_24u_0_7_7), 
           .COUT(co_mult_24u_24u_0_7_8), .S0(s_mult_24u_24u_0_7_25), .S1(s_mult_24u_24u_0_7_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_9 (.A0(s_mult_24u_24u_0_2_27), .A1(s_mult_24u_24u_0_2_28), 
           .B0(s_mult_24u_24u_0_3_27), .B1(s_mult_24u_24u_0_3_28), .CI(co_mult_24u_24u_0_7_8), 
           .COUT(co_mult_24u_24u_0_7_9), .S0(s_mult_24u_24u_0_7_27), .S1(s_mult_24u_24u_0_7_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_10 (.A0(s_mult_24u_24u_0_2_29), .A1(s_mult_24u_24u_0_2_30), 
           .B0(s_mult_24u_24u_0_3_29), .B1(s_mult_24u_24u_0_3_30), .CI(co_mult_24u_24u_0_7_9), 
           .COUT(co_mult_24u_24u_0_7_10), .S0(s_mult_24u_24u_0_7_29), .S1(s_mult_24u_24u_0_7_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_11 (.A0(s_mult_24u_24u_0_2_31), .A1(s_mult_24u_24u_0_2_32), 
           .B0(s_mult_24u_24u_0_3_31), .B1(s_mult_24u_24u_0_3_32), .CI(co_mult_24u_24u_0_7_10), 
           .COUT(co_mult_24u_24u_0_7_11), .S0(s_mult_24u_24u_0_7_31), .S1(s_mult_24u_24u_0_7_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_12 (.A0(s_mult_24u_24u_0_2_33), .A1(s_mult_24u_24u_0_2_34), 
           .B0(s_mult_24u_24u_0_3_33), .B1(s_mult_24u_24u_0_3_34), .CI(co_mult_24u_24u_0_7_11), 
           .COUT(co_mult_24u_24u_0_7_12), .S0(s_mult_24u_24u_0_7_33), .S1(s_mult_24u_24u_0_7_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_13 (.A0(s_mult_24u_24u_0_2_35), .A1(s_mult_24u_24u_0_2_36), 
           .B0(s_mult_24u_24u_0_3_35), .B1(s_mult_24u_24u_0_3_36), .CI(co_mult_24u_24u_0_7_12), 
           .COUT(co_mult_24u_24u_0_7_13), .S0(s_mult_24u_24u_0_7_35), .S1(s_mult_24u_24u_0_7_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_14 (.A0(s_mult_24u_24u_0_2_37), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_3_37), .B1(s_mult_24u_24u_0_3_38), .CI(co_mult_24u_24u_0_7_13), 
           .COUT(co_mult_24u_24u_0_7_14), .S0(s_mult_24u_24u_0_7_37), .S1(s_mult_24u_24u_0_7_38)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_3_39), .B1(s_mult_24u_24u_0_3_40), .CI(co_mult_24u_24u_0_7_14), 
           .COUT(co_mult_24u_24u_0_7_15), .S0(s_mult_24u_24u_0_7_39), .S1(s_mult_24u_24u_0_7_40)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_7_16 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_3_41), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_7_15), 
           .COUT(co_mult_24u_24u_0_7_16), .S0(s_mult_24u_24u_0_7_41), .S1(s_mult_24u_24u_0_7_42)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_7_17 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_7_16), 
           .S0(s_mult_24u_24u_0_7_43)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_8_1 (.A0(inputNumber[31]), .A1(s_mult_24u_24u_0_4_20), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_10_20), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_8_1), .S1(s_mult_24u_24u_0_8_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_2 (.A0(s_mult_24u_24u_0_4_21), .A1(s_mult_24u_24u_0_4_22), 
           .B0(mult_24u_24u_0_pp_10_21), .B1(s_mult_24u_24u_0_5_22), .CI(co_mult_24u_24u_0_8_1), 
           .COUT(co_mult_24u_24u_0_8_2), .S0(s_mult_24u_24u_0_8_21), .S1(s_mult_24u_24u_0_8_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_3 (.A0(s_mult_24u_24u_0_4_23), .A1(s_mult_24u_24u_0_4_24), 
           .B0(s_mult_24u_24u_0_5_23), .B1(s_mult_24u_24u_0_5_24), .CI(co_mult_24u_24u_0_8_2), 
           .COUT(co_mult_24u_24u_0_8_3), .S0(s_mult_24u_24u_0_8_23), .S1(s_mult_24u_24u_0_8_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_4 (.A0(s_mult_24u_24u_0_4_25), .A1(s_mult_24u_24u_0_4_26), 
           .B0(s_mult_24u_24u_0_5_25), .B1(s_mult_24u_24u_0_5_26), .CI(co_mult_24u_24u_0_8_3), 
           .COUT(co_mult_24u_24u_0_8_4), .S0(s_mult_24u_24u_0_8_25), .S1(s_mult_24u_24u_0_8_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_5 (.A0(s_mult_24u_24u_0_4_27), .A1(s_mult_24u_24u_0_4_28), 
           .B0(s_mult_24u_24u_0_5_27), .B1(s_mult_24u_24u_0_5_28), .CI(co_mult_24u_24u_0_8_4), 
           .COUT(co_mult_24u_24u_0_8_5), .S0(s_mult_24u_24u_0_8_27), .S1(s_mult_24u_24u_0_8_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_6 (.A0(s_mult_24u_24u_0_4_29), .A1(s_mult_24u_24u_0_4_30), 
           .B0(s_mult_24u_24u_0_5_29), .B1(s_mult_24u_24u_0_5_30), .CI(co_mult_24u_24u_0_8_5), 
           .COUT(co_mult_24u_24u_0_8_6), .S0(s_mult_24u_24u_0_8_29), .S1(s_mult_24u_24u_0_8_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_7 (.A0(s_mult_24u_24u_0_4_31), .A1(s_mult_24u_24u_0_4_32), 
           .B0(s_mult_24u_24u_0_5_31), .B1(s_mult_24u_24u_0_5_32), .CI(co_mult_24u_24u_0_8_6), 
           .COUT(co_mult_24u_24u_0_8_7), .S0(s_mult_24u_24u_0_8_31), .S1(s_mult_24u_24u_0_8_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_8 (.A0(s_mult_24u_24u_0_4_33), .A1(s_mult_24u_24u_0_4_34), 
           .B0(s_mult_24u_24u_0_5_33), .B1(s_mult_24u_24u_0_5_34), .CI(co_mult_24u_24u_0_8_7), 
           .COUT(co_mult_24u_24u_0_8_8), .S0(s_mult_24u_24u_0_8_33), .S1(s_mult_24u_24u_0_8_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_9 (.A0(s_mult_24u_24u_0_4_35), .A1(s_mult_24u_24u_0_4_36), 
           .B0(s_mult_24u_24u_0_5_35), .B1(s_mult_24u_24u_0_5_36), .CI(co_mult_24u_24u_0_8_8), 
           .COUT(co_mult_24u_24u_0_8_9), .S0(s_mult_24u_24u_0_8_35), .S1(s_mult_24u_24u_0_8_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_10 (.A0(s_mult_24u_24u_0_4_37), .A1(s_mult_24u_24u_0_4_38), 
           .B0(s_mult_24u_24u_0_5_37), .B1(s_mult_24u_24u_0_5_38), .CI(co_mult_24u_24u_0_8_9), 
           .COUT(co_mult_24u_24u_0_8_10), .S0(s_mult_24u_24u_0_8_37), .S1(s_mult_24u_24u_0_8_38)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_11 (.A0(s_mult_24u_24u_0_4_39), .A1(s_mult_24u_24u_0_4_40), 
           .B0(s_mult_24u_24u_0_5_39), .B1(s_mult_24u_24u_0_5_40), .CI(co_mult_24u_24u_0_8_10), 
           .COUT(co_mult_24u_24u_0_8_11), .S0(s_mult_24u_24u_0_8_39), .S1(s_mult_24u_24u_0_8_40)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_12 (.A0(s_mult_24u_24u_0_4_41), .A1(s_mult_24u_24u_0_4_42), 
           .B0(s_mult_24u_24u_0_5_41), .B1(s_mult_24u_24u_0_5_42), .CI(co_mult_24u_24u_0_8_11), 
           .COUT(co_mult_24u_24u_0_8_12), .S0(s_mult_24u_24u_0_8_41), .S1(s_mult_24u_24u_0_8_42)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_13 (.A0(s_mult_24u_24u_0_4_43), .A1(s_mult_24u_24u_0_4_44), 
           .B0(s_mult_24u_24u_0_5_43), .B1(s_mult_24u_24u_0_5_44), .CI(co_mult_24u_24u_0_8_12), 
           .COUT(co_mult_24u_24u_0_8_13), .S0(s_mult_24u_24u_0_8_43), .S1(s_mult_24u_24u_0_8_44)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_14 (.A0(s_mult_24u_24u_0_4_45), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_5_45), .B1(s_mult_24u_24u_0_5_46), .CI(co_mult_24u_24u_0_8_13), 
           .COUT(co_mult_24u_24u_0_8_14), .S0(s_mult_24u_24u_0_8_45), .S1(s_mult_24u_24u_0_8_46)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_8_15 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_5_47), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_8_14), 
           .S0(s_mult_24u_24u_0_8_47)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_9_1 (.A0(inputNumber[31]), .A1(s_mult_24u_24u_0_6_8), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_4_8), .CI(inputNumber[31]), 
           .COUT(co_mult_24u_24u_0_9_1)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_2 (.A0(s_mult_24u_24u_0_6_9), .A1(s_mult_24u_24u_0_6_10), 
           .B0(mult_24u_24u_0_pp_4_9), .B1(s_mult_24u_24u_0_2_10), .CI(co_mult_24u_24u_0_9_1), 
           .COUT(co_mult_24u_24u_0_9_2)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_3 (.A0(s_mult_24u_24u_0_6_11), .A1(s_mult_24u_24u_0_6_12), 
           .B0(s_mult_24u_24u_0_2_11), .B1(s_mult_24u_24u_0_7_12), .CI(co_mult_24u_24u_0_9_2), 
           .COUT(co_mult_24u_24u_0_9_3)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_4 (.A0(s_mult_24u_24u_0_6_13), .A1(s_mult_24u_24u_0_6_14), 
           .B0(s_mult_24u_24u_0_7_13), .B1(s_mult_24u_24u_0_7_14), .CI(co_mult_24u_24u_0_9_3), 
           .COUT(co_mult_24u_24u_0_9_4)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_5 (.A0(s_mult_24u_24u_0_6_15), .A1(s_mult_24u_24u_0_6_16), 
           .B0(s_mult_24u_24u_0_7_15), .B1(s_mult_24u_24u_0_7_16), .CI(co_mult_24u_24u_0_9_4), 
           .COUT(co_mult_24u_24u_0_9_5), .S1(s_mult_24u_24u_0_9_16)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_6 (.A0(s_mult_24u_24u_0_6_17), .A1(s_mult_24u_24u_0_6_18), 
           .B0(s_mult_24u_24u_0_7_17), .B1(s_mult_24u_24u_0_7_18), .CI(co_mult_24u_24u_0_9_5), 
           .COUT(co_mult_24u_24u_0_9_6), .S0(s_mult_24u_24u_0_9_17), .S1(s_mult_24u_24u_0_9_18)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_7 (.A0(s_mult_24u_24u_0_6_19), .A1(s_mult_24u_24u_0_6_20), 
           .B0(s_mult_24u_24u_0_7_19), .B1(s_mult_24u_24u_0_7_20), .CI(co_mult_24u_24u_0_9_6), 
           .COUT(co_mult_24u_24u_0_9_7), .S0(s_mult_24u_24u_0_9_19), .S1(s_mult_24u_24u_0_9_20)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_8 (.A0(s_mult_24u_24u_0_6_21), .A1(s_mult_24u_24u_0_6_22), 
           .B0(s_mult_24u_24u_0_7_21), .B1(s_mult_24u_24u_0_7_22), .CI(co_mult_24u_24u_0_9_7), 
           .COUT(co_mult_24u_24u_0_9_8), .S0(s_mult_24u_24u_0_9_21), .S1(s_mult_24u_24u_0_9_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_9 (.A0(s_mult_24u_24u_0_6_23), .A1(s_mult_24u_24u_0_6_24), 
           .B0(s_mult_24u_24u_0_7_23), .B1(s_mult_24u_24u_0_7_24), .CI(co_mult_24u_24u_0_9_8), 
           .COUT(co_mult_24u_24u_0_9_9), .S0(s_mult_24u_24u_0_9_23), .S1(s_mult_24u_24u_0_9_24)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_10 (.A0(s_mult_24u_24u_0_6_25), .A1(s_mult_24u_24u_0_6_26), 
           .B0(s_mult_24u_24u_0_7_25), .B1(s_mult_24u_24u_0_7_26), .CI(co_mult_24u_24u_0_9_9), 
           .COUT(co_mult_24u_24u_0_9_10), .S0(s_mult_24u_24u_0_9_25), .S1(s_mult_24u_24u_0_9_26)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_11 (.A0(s_mult_24u_24u_0_6_27), .A1(s_mult_24u_24u_0_6_28), 
           .B0(s_mult_24u_24u_0_7_27), .B1(s_mult_24u_24u_0_7_28), .CI(co_mult_24u_24u_0_9_10), 
           .COUT(co_mult_24u_24u_0_9_11), .S0(s_mult_24u_24u_0_9_27), .S1(s_mult_24u_24u_0_9_28)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_12 (.A0(s_mult_24u_24u_0_6_29), .A1(s_mult_24u_24u_0_6_30), 
           .B0(s_mult_24u_24u_0_7_29), .B1(s_mult_24u_24u_0_7_30), .CI(co_mult_24u_24u_0_9_11), 
           .COUT(co_mult_24u_24u_0_9_12), .S0(s_mult_24u_24u_0_9_29), .S1(s_mult_24u_24u_0_9_30)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_13 (.A0(s_mult_24u_24u_0_6_31), .A1(s_mult_24u_24u_0_6_32), 
           .B0(s_mult_24u_24u_0_7_31), .B1(s_mult_24u_24u_0_7_32), .CI(co_mult_24u_24u_0_9_12), 
           .COUT(co_mult_24u_24u_0_9_13), .S0(s_mult_24u_24u_0_9_31), .S1(s_mult_24u_24u_0_9_32)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_14 (.A0(s_mult_24u_24u_0_6_33), .A1(s_mult_24u_24u_0_6_34), 
           .B0(s_mult_24u_24u_0_7_33), .B1(s_mult_24u_24u_0_7_34), .CI(co_mult_24u_24u_0_9_13), 
           .COUT(co_mult_24u_24u_0_9_14), .S0(s_mult_24u_24u_0_9_33), .S1(s_mult_24u_24u_0_9_34)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_15 (.A0(s_mult_24u_24u_0_6_35), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_7_35), .B1(s_mult_24u_24u_0_7_36), .CI(co_mult_24u_24u_0_9_14), 
           .COUT(co_mult_24u_24u_0_9_15), .S0(s_mult_24u_24u_0_9_35), .S1(s_mult_24u_24u_0_9_36)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_16 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_7_37), .B1(s_mult_24u_24u_0_7_38), .CI(co_mult_24u_24u_0_9_15), 
           .COUT(co_mult_24u_24u_0_9_16), .S0(s_mult_24u_24u_0_9_37), .S1(s_mult_24u_24u_0_9_38)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_17 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_7_39), .B1(s_mult_24u_24u_0_7_40), .CI(co_mult_24u_24u_0_9_16), 
           .COUT(co_mult_24u_24u_0_9_17), .S0(s_mult_24u_24u_0_9_39), .S1(s_mult_24u_24u_0_9_40)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_18 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_7_41), .B1(s_mult_24u_24u_0_7_42), .CI(co_mult_24u_24u_0_9_17), 
           .COUT(co_mult_24u_24u_0_9_18), .S0(s_mult_24u_24u_0_9_41), .S1(s_mult_24u_24u_0_9_42)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_add_9_19 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_7_43), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_9_18), 
           .COUT(co_mult_24u_24u_0_9_19), .S0(s_mult_24u_24u_0_9_43), .S1(s_mult_24u_24u_0_9_44)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_mult_24u_24u_0_9_20 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(co_mult_24u_24u_0_9_19), 
           .S0(s_mult_24u_24u_0_9_45)) /* synthesis syn_instantiated=1 */ ;
    FADD2B Cadd_t_mult_24u_24u_0_10_1 (.A0(inputNumber[31]), .A1(s_mult_24u_24u_0_9_16), 
           .B0(inputNumber[31]), .B1(mult_24u_24u_0_pp_8_16), .CI(inputNumber[31]), 
           .COUT(co_t_mult_24u_24u_0_10_1)) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_2 (.A0(s_mult_24u_24u_0_9_17), .A1(s_mult_24u_24u_0_9_18), 
           .B0(mult_24u_24u_0_pp_8_17), .B1(s_mult_24u_24u_0_4_18), .CI(co_t_mult_24u_24u_0_10_1), 
           .COUT(co_t_mult_24u_24u_0_10_2)) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_3 (.A0(s_mult_24u_24u_0_9_19), .A1(s_mult_24u_24u_0_9_20), 
           .B0(s_mult_24u_24u_0_4_19), .B1(s_mult_24u_24u_0_8_20), .CI(co_t_mult_24u_24u_0_10_2), 
           .COUT(co_t_mult_24u_24u_0_10_3)) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_4 (.A0(s_mult_24u_24u_0_9_21), .A1(s_mult_24u_24u_0_9_22), 
           .B0(s_mult_24u_24u_0_8_21), .B1(s_mult_24u_24u_0_8_22), .CI(co_t_mult_24u_24u_0_10_3), 
           .COUT(co_t_mult_24u_24u_0_10_4), .S0(prod[21]), .S1(prod[22])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_5 (.A0(s_mult_24u_24u_0_9_23), .A1(s_mult_24u_24u_0_9_24), 
           .B0(s_mult_24u_24u_0_8_23), .B1(s_mult_24u_24u_0_8_24), .CI(co_t_mult_24u_24u_0_10_4), 
           .COUT(co_t_mult_24u_24u_0_10_5), .S0(prod[23]), .S1(prod[24])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_6 (.A0(s_mult_24u_24u_0_9_25), .A1(s_mult_24u_24u_0_9_26), 
           .B0(s_mult_24u_24u_0_8_25), .B1(s_mult_24u_24u_0_8_26), .CI(co_t_mult_24u_24u_0_10_5), 
           .COUT(co_t_mult_24u_24u_0_10_6), .S0(prod[25]), .S1(prod[26])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_7 (.A0(s_mult_24u_24u_0_9_27), .A1(s_mult_24u_24u_0_9_28), 
           .B0(s_mult_24u_24u_0_8_27), .B1(s_mult_24u_24u_0_8_28), .CI(co_t_mult_24u_24u_0_10_6), 
           .COUT(co_t_mult_24u_24u_0_10_7), .S0(prod[27]), .S1(prod[28])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_8 (.A0(s_mult_24u_24u_0_9_29), .A1(s_mult_24u_24u_0_9_30), 
           .B0(s_mult_24u_24u_0_8_29), .B1(s_mult_24u_24u_0_8_30), .CI(co_t_mult_24u_24u_0_10_7), 
           .COUT(co_t_mult_24u_24u_0_10_8), .S0(prod[29]), .S1(prod[30])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_9 (.A0(s_mult_24u_24u_0_9_31), .A1(s_mult_24u_24u_0_9_32), 
           .B0(s_mult_24u_24u_0_8_31), .B1(s_mult_24u_24u_0_8_32), .CI(co_t_mult_24u_24u_0_10_8), 
           .COUT(co_t_mult_24u_24u_0_10_9), .S0(prod[31]), .S1(prod[32])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_10 (.A0(s_mult_24u_24u_0_9_33), .A1(s_mult_24u_24u_0_9_34), 
           .B0(s_mult_24u_24u_0_8_33), .B1(s_mult_24u_24u_0_8_34), .CI(co_t_mult_24u_24u_0_10_9), 
           .COUT(co_t_mult_24u_24u_0_10_10), .S0(prod[33]), .S1(prod[34])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_11 (.A0(s_mult_24u_24u_0_9_35), .A1(s_mult_24u_24u_0_9_36), 
           .B0(s_mult_24u_24u_0_8_35), .B1(s_mult_24u_24u_0_8_36), .CI(co_t_mult_24u_24u_0_10_10), 
           .COUT(co_t_mult_24u_24u_0_10_11), .S0(prod[35]), .S1(prod[36])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_12 (.A0(s_mult_24u_24u_0_9_37), .A1(s_mult_24u_24u_0_9_38), 
           .B0(s_mult_24u_24u_0_8_37), .B1(s_mult_24u_24u_0_8_38), .CI(co_t_mult_24u_24u_0_10_11), 
           .COUT(co_t_mult_24u_24u_0_10_12), .S0(prod[37]), .S1(prod[38])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_13 (.A0(s_mult_24u_24u_0_9_39), .A1(s_mult_24u_24u_0_9_40), 
           .B0(s_mult_24u_24u_0_8_39), .B1(s_mult_24u_24u_0_8_40), .CI(co_t_mult_24u_24u_0_10_12), 
           .COUT(co_t_mult_24u_24u_0_10_13), .S0(prod[39]), .S1(prod[40])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_14 (.A0(s_mult_24u_24u_0_9_41), .A1(s_mult_24u_24u_0_9_42), 
           .B0(s_mult_24u_24u_0_8_41), .B1(s_mult_24u_24u_0_8_42), .CI(co_t_mult_24u_24u_0_10_13), 
           .COUT(co_t_mult_24u_24u_0_10_14), .S0(prod[41]), .S1(prod[42])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_15 (.A0(s_mult_24u_24u_0_9_43), .A1(s_mult_24u_24u_0_9_44), 
           .B0(s_mult_24u_24u_0_8_43), .B1(s_mult_24u_24u_0_8_44), .CI(co_t_mult_24u_24u_0_10_14), 
           .COUT(co_t_mult_24u_24u_0_10_15), .S0(prod[43]), .S1(prod[44])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_16 (.A0(s_mult_24u_24u_0_9_45), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_8_45), .B1(s_mult_24u_24u_0_8_46), .CI(co_t_mult_24u_24u_0_10_15), 
           .COUT(co_t_mult_24u_24u_0_10_16), .S0(prod[45]), .S1(prod[46])) /* synthesis syn_instantiated=1 */ ;
    FADD2B t_mult_24u_24u_0_add_10_17 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(s_mult_24u_24u_0_8_47), .B1(inputNumber[31]), .CI(co_t_mult_24u_24u_0_10_16), 
           .S0(prod[47])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mult_24u_24u_0_cin_lr_0), .CO(mco), .P1(mult_24u_24u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco), .CO(mco_1), .P0(mult_24u_24u_0_pp_0_3), .P1(mult_24u_24u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_1), .CO(mco_2), .P0(mult_24u_24u_0_pp_0_5), .P1(mult_24u_24u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_2), .CO(mco_3), .P0(mult_24u_24u_0_pp_0_7), .P1(mult_24u_24u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_3), .CO(mco_4), .P0(mult_24u_24u_0_pp_0_9), .P1(mult_24u_24u_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_4), .CO(mco_5), .P0(mult_24u_24u_0_pp_0_11), .P1(mult_24u_24u_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_5), .CO(mco_6), .P0(mult_24u_24u_0_pp_0_13), .P1(mult_24u_24u_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_6), .CO(mco_7), .P0(mult_24u_24u_0_pp_0_15), .P1(mult_24u_24u_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_7), .CO(mco_8), .P0(mult_24u_24u_0_pp_0_17), .P1(mult_24u_24u_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_8), .CO(mco_9), .P0(mult_24u_24u_0_pp_0_19), .P1(mult_24u_24u_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_9), .CO(mco_10), .P0(mult_24u_24u_0_pp_0_21), .P1(mult_24u_24u_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_0_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[1]), 
          .B1(B_int_adj_725[0]), .B2(B_int_adj_725[1]), .B3(B_int_adj_725[0]), 
          .CI(mco_10), .CO(mfco), .P0(mult_24u_24u_0_pp_0_23), .P1(mult_24u_24u_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mult_24u_24u_0_cin_lr_2), .CO(mco_11), .P0(mult_24u_24u_0_pp_1_3), 
          .P1(mult_24u_24u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_11), .CO(mco_12), .P0(mult_24u_24u_0_pp_1_5), .P1(mult_24u_24u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_12), .CO(mco_13), .P0(mult_24u_24u_0_pp_1_7), .P1(mult_24u_24u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_13), .CO(mco_14), .P0(mult_24u_24u_0_pp_1_9), .P1(mult_24u_24u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_14), .CO(mco_15), .P0(mult_24u_24u_0_pp_1_11), .P1(mult_24u_24u_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_15), .CO(mco_16), .P0(mult_24u_24u_0_pp_1_13), .P1(mult_24u_24u_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_16), .CO(mco_17), .P0(mult_24u_24u_0_pp_1_15), .P1(mult_24u_24u_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_17), .CO(mco_18), .P0(mult_24u_24u_0_pp_1_17), .P1(mult_24u_24u_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_18), .CO(mco_19), .P0(mult_24u_24u_0_pp_1_19), .P1(mult_24u_24u_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_19), .CO(mco_20), .P0(mult_24u_24u_0_pp_1_21), .P1(mult_24u_24u_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_20), .CO(mco_21), .P0(mult_24u_24u_0_pp_1_23), .P1(mult_24u_24u_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_2_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[3]), 
          .B1(B_int_adj_725[2]), .B2(B_int_adj_725[3]), .B3(B_int_adj_725[2]), 
          .CI(mco_21), .CO(mfco_1), .P0(mult_24u_24u_0_pp_1_25), .P1(mult_24u_24u_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mult_24u_24u_0_cin_lr_4), .CO(mco_22), .P0(mult_24u_24u_0_pp_2_5), 
          .P1(mult_24u_24u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_22), .CO(mco_23), .P0(mult_24u_24u_0_pp_2_7), .P1(mult_24u_24u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_23), .CO(mco_24), .P0(mult_24u_24u_0_pp_2_9), .P1(mult_24u_24u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_24), .CO(mco_25), .P0(mult_24u_24u_0_pp_2_11), .P1(mult_24u_24u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_25), .CO(mco_26), .P0(mult_24u_24u_0_pp_2_13), .P1(mult_24u_24u_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_26), .CO(mco_27), .P0(mult_24u_24u_0_pp_2_15), .P1(mult_24u_24u_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_27), .CO(mco_28), .P0(mult_24u_24u_0_pp_2_17), .P1(mult_24u_24u_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_28), .CO(mco_29), .P0(mult_24u_24u_0_pp_2_19), .P1(mult_24u_24u_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_29), .CO(mco_30), .P0(mult_24u_24u_0_pp_2_21), .P1(mult_24u_24u_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_30), .CO(mco_31), .P0(mult_24u_24u_0_pp_2_23), .P1(mult_24u_24u_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_31), .CO(mco_32), .P0(mult_24u_24u_0_pp_2_25), .P1(mult_24u_24u_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_4_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[5]), 
          .B1(B_int_adj_725[4]), .B2(B_int_adj_725[5]), .B3(B_int_adj_725[4]), 
          .CI(mco_32), .CO(mfco_2), .P0(mult_24u_24u_0_pp_2_27), .P1(mult_24u_24u_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mult_24u_24u_0_cin_lr_6), .CO(mco_33), .P0(mult_24u_24u_0_pp_3_7), 
          .P1(mult_24u_24u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_33), .CO(mco_34), .P0(mult_24u_24u_0_pp_3_9), .P1(mult_24u_24u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_34), .CO(mco_35), .P0(mult_24u_24u_0_pp_3_11), .P1(mult_24u_24u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_35), .CO(mco_36), .P0(mult_24u_24u_0_pp_3_13), .P1(mult_24u_24u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_36), .CO(mco_37), .P0(mult_24u_24u_0_pp_3_15), .P1(mult_24u_24u_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_37), .CO(mco_38), .P0(mult_24u_24u_0_pp_3_17), .P1(mult_24u_24u_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_38), .CO(mco_39), .P0(mult_24u_24u_0_pp_3_19), .P1(mult_24u_24u_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_39), .CO(mco_40), .P0(mult_24u_24u_0_pp_3_21), .P1(mult_24u_24u_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_40), .CO(mco_41), .P0(mult_24u_24u_0_pp_3_23), .P1(mult_24u_24u_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_41), .CO(mco_42), .P0(mult_24u_24u_0_pp_3_25), .P1(mult_24u_24u_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_42), .CO(mco_43), .P0(mult_24u_24u_0_pp_3_27), .P1(mult_24u_24u_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_6_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[7]), 
          .B1(B_int_adj_725[6]), .B2(B_int_adj_725[7]), .B3(B_int_adj_725[6]), 
          .CI(mco_43), .CO(mfco_3), .P0(mult_24u_24u_0_pp_3_29), .P1(mult_24u_24u_0_pp_3_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mult_24u_24u_0_cin_lr_8), .CO(mco_44), .P0(mult_24u_24u_0_pp_4_9), 
          .P1(mult_24u_24u_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_44), .CO(mco_45), .P0(mult_24u_24u_0_pp_4_11), .P1(mult_24u_24u_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_45), .CO(mco_46), .P0(mult_24u_24u_0_pp_4_13), .P1(mult_24u_24u_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_46), .CO(mco_47), .P0(mult_24u_24u_0_pp_4_15), .P1(mult_24u_24u_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_47), .CO(mco_48), .P0(mult_24u_24u_0_pp_4_17), .P1(mult_24u_24u_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_48), .CO(mco_49), .P0(mult_24u_24u_0_pp_4_19), .P1(mult_24u_24u_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_49), .CO(mco_50), .P0(mult_24u_24u_0_pp_4_21), .P1(mult_24u_24u_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_50), .CO(mco_51), .P0(mult_24u_24u_0_pp_4_23), .P1(mult_24u_24u_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_51), .CO(mco_52), .P0(mult_24u_24u_0_pp_4_25), .P1(mult_24u_24u_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_52), .CO(mco_53), .P0(mult_24u_24u_0_pp_4_27), .P1(mult_24u_24u_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_53), .CO(mco_54), .P0(mult_24u_24u_0_pp_4_29), .P1(mult_24u_24u_0_pp_4_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_8_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[9]), 
          .B1(B_int_adj_725[8]), .B2(B_int_adj_725[9]), .B3(B_int_adj_725[8]), 
          .CI(mco_54), .CO(mfco_4), .P0(mult_24u_24u_0_pp_4_31), .P1(mult_24u_24u_0_pp_4_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mult_24u_24u_0_cin_lr_10), .CO(mco_55), .P0(mult_24u_24u_0_pp_5_11), 
          .P1(mult_24u_24u_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_55), .CO(mco_56), .P0(mult_24u_24u_0_pp_5_13), .P1(mult_24u_24u_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_56), .CO(mco_57), .P0(mult_24u_24u_0_pp_5_15), .P1(mult_24u_24u_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_57), .CO(mco_58), .P0(mult_24u_24u_0_pp_5_17), .P1(mult_24u_24u_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_58), .CO(mco_59), .P0(mult_24u_24u_0_pp_5_19), .P1(mult_24u_24u_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_59), .CO(mco_60), .P0(mult_24u_24u_0_pp_5_21), .P1(mult_24u_24u_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_60), .CO(mco_61), .P0(mult_24u_24u_0_pp_5_23), .P1(mult_24u_24u_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_61), .CO(mco_62), .P0(mult_24u_24u_0_pp_5_25), .P1(mult_24u_24u_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_62), .CO(mco_63), .P0(mult_24u_24u_0_pp_5_27), .P1(mult_24u_24u_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_63), .CO(mco_64), .P0(mult_24u_24u_0_pp_5_29), .P1(mult_24u_24u_0_pp_5_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_64), .CO(mco_65), .P0(mult_24u_24u_0_pp_5_31), .P1(mult_24u_24u_0_pp_5_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_10_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[11]), 
          .B1(B_int_adj_725[10]), .B2(B_int_adj_725[11]), .B3(B_int_adj_725[10]), 
          .CI(mco_65), .CO(mfco_5), .P0(mult_24u_24u_0_pp_5_33), .P1(mult_24u_24u_0_pp_5_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mult_24u_24u_0_cin_lr_12), .CO(mco_66), .P0(mult_24u_24u_0_pp_6_13), 
          .P1(mult_24u_24u_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_66), .CO(mco_67), .P0(mult_24u_24u_0_pp_6_15), .P1(mult_24u_24u_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_67), .CO(mco_68), .P0(mult_24u_24u_0_pp_6_17), .P1(mult_24u_24u_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_68), .CO(mco_69), .P0(mult_24u_24u_0_pp_6_19), .P1(mult_24u_24u_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_69), .CO(mco_70), .P0(mult_24u_24u_0_pp_6_21), .P1(mult_24u_24u_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_70), .CO(mco_71), .P0(mult_24u_24u_0_pp_6_23), .P1(mult_24u_24u_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_71), .CO(mco_72), .P0(mult_24u_24u_0_pp_6_25), .P1(mult_24u_24u_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_72), .CO(mco_73), .P0(mult_24u_24u_0_pp_6_27), .P1(mult_24u_24u_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_73), .CO(mco_74), .P0(mult_24u_24u_0_pp_6_29), .P1(mult_24u_24u_0_pp_6_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_74), .CO(mco_75), .P0(mult_24u_24u_0_pp_6_31), .P1(mult_24u_24u_0_pp_6_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_75), .CO(mco_76), .P0(mult_24u_24u_0_pp_6_33), .P1(mult_24u_24u_0_pp_6_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_12_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[13]), 
          .B1(B_int_adj_725[12]), .B2(B_int_adj_725[13]), .B3(B_int_adj_725[12]), 
          .CI(mco_76), .CO(mfco_6), .P0(mult_24u_24u_0_pp_6_35), .P1(mult_24u_24u_0_pp_6_36)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mult_24u_24u_0_cin_lr_14), .CO(mco_77), .P0(mult_24u_24u_0_pp_7_15), 
          .P1(mult_24u_24u_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_77), .CO(mco_78), .P0(mult_24u_24u_0_pp_7_17), .P1(mult_24u_24u_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_78), .CO(mco_79), .P0(mult_24u_24u_0_pp_7_19), .P1(mult_24u_24u_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_79), .CO(mco_80), .P0(mult_24u_24u_0_pp_7_21), .P1(mult_24u_24u_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_80), .CO(mco_81), .P0(mult_24u_24u_0_pp_7_23), .P1(mult_24u_24u_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_81), .CO(mco_82), .P0(mult_24u_24u_0_pp_7_25), .P1(mult_24u_24u_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_82), .CO(mco_83), .P0(mult_24u_24u_0_pp_7_27), .P1(mult_24u_24u_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_83), .CO(mco_84), .P0(mult_24u_24u_0_pp_7_29), .P1(mult_24u_24u_0_pp_7_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_84), .CO(mco_85), .P0(mult_24u_24u_0_pp_7_31), .P1(mult_24u_24u_0_pp_7_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_85), .CO(mco_86), .P0(mult_24u_24u_0_pp_7_33), .P1(mult_24u_24u_0_pp_7_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_86), .CO(mco_87), .P0(mult_24u_24u_0_pp_7_35), .P1(mult_24u_24u_0_pp_7_36)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_14_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[15]), 
          .B1(B_int_adj_725[14]), .B2(B_int_adj_725[15]), .B3(B_int_adj_725[14]), 
          .CI(mco_87), .CO(mfco_7), .P0(mult_24u_24u_0_pp_7_37), .P1(mult_24u_24u_0_pp_7_38)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mult_24u_24u_0_cin_lr_16), .CO(mco_88), .P0(mult_24u_24u_0_pp_8_17), 
          .P1(mult_24u_24u_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_88), .CO(mco_89), .P0(mult_24u_24u_0_pp_8_19), .P1(mult_24u_24u_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_89), .CO(mco_90), .P0(mult_24u_24u_0_pp_8_21), .P1(mult_24u_24u_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_90), .CO(mco_91), .P0(mult_24u_24u_0_pp_8_23), .P1(mult_24u_24u_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_91), .CO(mco_92), .P0(mult_24u_24u_0_pp_8_25), .P1(mult_24u_24u_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_92), .CO(mco_93), .P0(mult_24u_24u_0_pp_8_27), .P1(mult_24u_24u_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_93), .CO(mco_94), .P0(mult_24u_24u_0_pp_8_29), .P1(mult_24u_24u_0_pp_8_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_94), .CO(mco_95), .P0(mult_24u_24u_0_pp_8_31), .P1(mult_24u_24u_0_pp_8_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_95), .CO(mco_96), .P0(mult_24u_24u_0_pp_8_33), .P1(mult_24u_24u_0_pp_8_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_96), .CO(mco_97), .P0(mult_24u_24u_0_pp_8_35), .P1(mult_24u_24u_0_pp_8_36)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_97), .CO(mco_98), .P0(mult_24u_24u_0_pp_8_37), .P1(mult_24u_24u_0_pp_8_38)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_16_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[17]), 
          .B1(B_int_adj_725[16]), .B2(B_int_adj_725[17]), .B3(B_int_adj_725[16]), 
          .CI(mco_98), .CO(mfco_8), .P0(mult_24u_24u_0_pp_8_39), .P1(mult_24u_24u_0_pp_8_40)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mult_24u_24u_0_cin_lr_18), .CO(mco_99), .P0(mult_24u_24u_0_pp_9_19), 
          .P1(mult_24u_24u_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_99), .CO(mco_100), .P0(mult_24u_24u_0_pp_9_21), .P1(mult_24u_24u_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_100), .CO(mco_101), .P0(mult_24u_24u_0_pp_9_23), .P1(mult_24u_24u_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_101), .CO(mco_102), .P0(mult_24u_24u_0_pp_9_25), .P1(mult_24u_24u_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_102), .CO(mco_103), .P0(mult_24u_24u_0_pp_9_27), .P1(mult_24u_24u_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_103), .CO(mco_104), .P0(mult_24u_24u_0_pp_9_29), .P1(mult_24u_24u_0_pp_9_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_104), .CO(mco_105), .P0(mult_24u_24u_0_pp_9_31), .P1(mult_24u_24u_0_pp_9_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_105), .CO(mco_106), .P0(mult_24u_24u_0_pp_9_33), .P1(mult_24u_24u_0_pp_9_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_106), .CO(mco_107), .P0(mult_24u_24u_0_pp_9_35), .P1(mult_24u_24u_0_pp_9_36)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_107), .CO(mco_108), .P0(mult_24u_24u_0_pp_9_37), .P1(mult_24u_24u_0_pp_9_38)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_108), .CO(mco_109), .P0(mult_24u_24u_0_pp_9_39), .P1(mult_24u_24u_0_pp_9_40)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_18_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[19]), 
          .B1(B_int_adj_725[18]), .B2(B_int_adj_725[19]), .B3(B_int_adj_725[18]), 
          .CI(mco_109), .CO(mfco_9), .P0(mult_24u_24u_0_pp_9_41), .P1(mult_24u_24u_0_pp_9_42)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mult_24u_24u_0_cin_lr_20), .CO(mco_110), .P0(mult_24u_24u_0_pp_10_21), 
          .P1(mult_24u_24u_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_110), .CO(mco_111), .P0(mult_24u_24u_0_pp_10_23), .P1(mult_24u_24u_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_111), .CO(mco_112), .P0(mult_24u_24u_0_pp_10_25), .P1(mult_24u_24u_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_112), .CO(mco_113), .P0(mult_24u_24u_0_pp_10_27), .P1(mult_24u_24u_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_113), .CO(mco_114), .P0(mult_24u_24u_0_pp_10_29), .P1(mult_24u_24u_0_pp_10_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_114), .CO(mco_115), .P0(mult_24u_24u_0_pp_10_31), .P1(mult_24u_24u_0_pp_10_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_115), .CO(mco_116), .P0(mult_24u_24u_0_pp_10_33), .P1(mult_24u_24u_0_pp_10_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_116), .CO(mco_117), .P0(mult_24u_24u_0_pp_10_35), .P1(mult_24u_24u_0_pp_10_36)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_117), .CO(mco_118), .P0(mult_24u_24u_0_pp_10_37), .P1(mult_24u_24u_0_pp_10_38)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_118), .CO(mco_119), .P0(mult_24u_24u_0_pp_10_39), .P1(mult_24u_24u_0_pp_10_40)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_119), .CO(mco_120), .P0(mult_24u_24u_0_pp_10_41), .P1(mult_24u_24u_0_pp_10_42)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_20_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(B_int_adj_725[21]), 
          .B1(B_int_adj_725[20]), .B2(B_int_adj_725[21]), .B3(B_int_adj_725[20]), 
          .CI(mco_120), .CO(mfco_10), .P0(mult_24u_24u_0_pp_10_43), .P1(mult_24u_24u_0_pp_10_44)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_0 (.A0(A_int_adj_724[0]), .A1(A_int_adj_724[1]), 
          .A2(A_int_adj_724[1]), .A3(A_int_adj_724[2]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mult_24u_24u_0_cin_lr_22), .CO(mco_121), .P0(mult_24u_24u_0_pp_11_23), 
          .P1(mult_24u_24u_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_1 (.A0(A_int_adj_724[2]), .A1(A_int_adj_724[3]), 
          .A2(A_int_adj_724[3]), .A3(A_int_adj_724[4]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_121), .CO(mco_122), .P0(mult_24u_24u_0_pp_11_25), .P1(mult_24u_24u_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_2 (.A0(A_int_adj_724[4]), .A1(A_int_adj_724[5]), 
          .A2(A_int_adj_724[5]), .A3(A_int_adj_724[6]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_122), .CO(mco_123), .P0(mult_24u_24u_0_pp_11_27), .P1(mult_24u_24u_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_3 (.A0(A_int_adj_724[6]), .A1(A_int_adj_724[7]), 
          .A2(A_int_adj_724[7]), .A3(A_int_adj_724[8]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_123), .CO(mco_124), .P0(mult_24u_24u_0_pp_11_29), .P1(mult_24u_24u_0_pp_11_30)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_4 (.A0(A_int_adj_724[8]), .A1(A_int_adj_724[9]), 
          .A2(A_int_adj_724[9]), .A3(A_int_adj_724[10]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_124), .CO(mco_125), .P0(mult_24u_24u_0_pp_11_31), .P1(mult_24u_24u_0_pp_11_32)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_5 (.A0(A_int_adj_724[10]), .A1(A_int_adj_724[11]), 
          .A2(A_int_adj_724[11]), .A3(A_int_adj_724[12]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_125), .CO(mco_126), .P0(mult_24u_24u_0_pp_11_33), .P1(mult_24u_24u_0_pp_11_34)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_6 (.A0(A_int_adj_724[12]), .A1(A_int_adj_724[13]), 
          .A2(A_int_adj_724[13]), .A3(A_int_adj_724[14]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_126), .CO(mco_127), .P0(mult_24u_24u_0_pp_11_35), .P1(mult_24u_24u_0_pp_11_36)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_7 (.A0(A_int_adj_724[14]), .A1(A_int_adj_724[15]), 
          .A2(A_int_adj_724[15]), .A3(A_int_adj_724[16]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_127), .CO(mco_128), .P0(mult_24u_24u_0_pp_11_37), .P1(mult_24u_24u_0_pp_11_38)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_8 (.A0(A_int_adj_724[16]), .A1(A_int_adj_724[17]), 
          .A2(A_int_adj_724[17]), .A3(A_int_adj_724[18]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_128), .CO(mco_129), .P0(mult_24u_24u_0_pp_11_39), .P1(mult_24u_24u_0_pp_11_40)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_9 (.A0(A_int_adj_724[18]), .A1(A_int_adj_724[19]), 
          .A2(A_int_adj_724[19]), .A3(A_int_adj_724[20]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_129), .CO(mco_130), .P0(mult_24u_24u_0_pp_11_41), .P1(mult_24u_24u_0_pp_11_42)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_10 (.A0(A_int_adj_724[20]), .A1(A_int_adj_724[21]), 
          .A2(A_int_adj_724[21]), .A3(A_int_adj_724[22]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_130), .CO(mco_131), .P0(mult_24u_24u_0_pp_11_43), .P1(mult_24u_24u_0_pp_11_44)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_24u_24u_0_mult_22_11 (.A0(A_int_adj_724[22]), .A1(inputNumber[2]), 
          .A2(inputNumber[2]), .A3(inputNumber[31]), .B0(inputNumber[2]), 
          .B1(B_int_adj_725[22]), .B2(inputNumber[2]), .B3(B_int_adj_725[22]), 
          .CI(mco_131), .CO(mfco_11), .P0(mult_24u_24u_0_pp_11_45), .P1(mult_24u_24u_0_pp_11_46)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t6 (.A(A_int_adj_724[0]), .B(B_int_adj_725[10]), .Z(mult_24u_24u_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t5 (.A(A_int_adj_724[0]), .B(B_int_adj_725[12]), .Z(mult_24u_24u_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t4 (.A(A_int_adj_724[0]), .B(B_int_adj_725[14]), .Z(mult_24u_24u_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t3 (.A(A_int_adj_724[0]), .B(B_int_adj_725[16]), .Z(mult_24u_24u_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t2 (.A(A_int_adj_724[0]), .B(B_int_adj_725[18]), .Z(mult_24u_24u_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t1 (.A(A_int_adj_724[0]), .B(B_int_adj_725[20]), .Z(mult_24u_24u_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;
    AND2 AND2_t0_adj_985 (.A(A_int_adj_724[0]), .B(B_int_adj_725[22]), .Z(mult_24u_24u_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_24u_24u_0_cin_lr_add_0 (.A0(inputNumber[31]), .A1(inputNumber[31]), 
           .B0(inputNumber[31]), .B1(inputNumber[31]), .CI(inputNumber[31]), 
           .COUT(mult_24u_24u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;
    LUT4 i12289_2_lut_4_lut (.A(n73809), .B(n1148[0]), .C(SDA_c), .D(n1148[5]), 
         .Z(n23979)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i12289_2_lut_4_lut.init = 16'h0200;
    LUT4 i55085_3_lut_rep_774 (.A(n73809), .B(n1148[0]), .C(SDA_c), .Z(n70744)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i55085_3_lut_rep_774.init = 16'h0202;
    AND2 AND2_t32 (.A(i[0]), .B(inputNumber[31]), .Z(n898[0])) /* synthesis syn_instantiated=1 */ ;
    IB SDA_pad (.I(SDA), .O(SDA_c));
    ND2 ND2_t30 (.A(i[0]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_0_n0)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t29 (.A(i[3]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_1_n1)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t28 (.A(i[2]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_1_n0)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t27 (.A(i[5]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_2_n1)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t26 (.A(i[4]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_2_n0)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t25 (.A(i[7]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_3_n1)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t24 (.A(i[6]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_3_n0)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t23 (.A(i[9]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_4_n1)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t22 (.A(i[8]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_4_n0)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t21 (.A(i[11]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_5_n1)) /* synthesis syn_instantiated=1 */ ;
    ND2 ND2_t20 (.A(i[10]), .B(n14049[1]), .Z(mult_32s_2s_0_mult_0_5_n0)) /* synthesis syn_instantiated=1 */ ;
    FADD2B mult_32s_2s_0_cin_lr_add (.A0(inputNumber[2]), .A1(inputNumber[2]), 
           .B0(inputNumber[2]), .B1(inputNumber[2]), .CI(inputNumber[31]), 
           .COUT(mult_32s_2s_0_cin_lr)) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_32s_2s_0_mult_0_0 (.A0(mult_32s_2s_0_mult_0_0_n0), .A1(i[1]), 
          .A2(mult_32s_2s_0_mult_0_0_n1), .A3(i[2]), .B0(inputNumber[2]), 
          .B1(inputNumber[31]), .B2(inputNumber[2]), .B3(inputNumber[31]), 
          .CI(mult_32s_2s_0_cin_lr), .CO(mco_adj_608), .P0(n898[1]), .P1(n898[2])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_32s_2s_0_mult_0_1 (.A0(mult_32s_2s_0_mult_0_1_n0), .A1(i[3]), 
          .A2(mult_32s_2s_0_mult_0_1_n1), .A3(i[4]), .B0(inputNumber[2]), 
          .B1(inputNumber[31]), .B2(inputNumber[2]), .B3(inputNumber[31]), 
          .CI(mco_adj_608), .CO(mco_1_adj_609), .P0(n898[3]), .P1(n898[4])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_32s_2s_0_mult_0_2 (.A0(mult_32s_2s_0_mult_0_2_n0), .A1(i[5]), 
          .A2(mult_32s_2s_0_mult_0_2_n1), .A3(i[6]), .B0(inputNumber[2]), 
          .B1(inputNumber[31]), .B2(inputNumber[2]), .B3(inputNumber[31]), 
          .CI(mco_1_adj_609), .CO(mco_2_adj_610), .P0(n898[5]), .P1(n898[6])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_32s_2s_0_mult_0_3 (.A0(mult_32s_2s_0_mult_0_3_n0), .A1(i[7]), 
          .A2(mult_32s_2s_0_mult_0_3_n1), .A3(i[8]), .B0(inputNumber[2]), 
          .B1(inputNumber[31]), .B2(inputNumber[2]), .B3(inputNumber[31]), 
          .CI(mco_2_adj_610), .CO(mco_3_adj_611), .P0(n898[7]), .P1(n898[8])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_32s_2s_0_mult_0_4 (.A0(mult_32s_2s_0_mult_0_4_n0), .A1(i[9]), 
          .A2(mult_32s_2s_0_mult_0_4_n1), .A3(i[10]), .B0(inputNumber[2]), 
          .B1(inputNumber[31]), .B2(inputNumber[2]), .B3(inputNumber[31]), 
          .CI(mco_3_adj_611), .CO(mco_4_adj_612), .P0(n898[9]), .P1(n898[10])) /* synthesis syn_instantiated=1 */ ;
    MULT2 mult_32s_2s_0_mult_0_5 (.A0(mult_32s_2s_0_mult_0_5_n0), .A1(i[11]), 
          .A2(mult_32s_2s_0_mult_0_5_n1), .A3(i[12]), .B0(inputNumber[2]), 
          .B1(inputNumber[31]), .B2(inputNumber[2]), .B3(inputNumber[31]), 
          .CI(mco_4_adj_612), .P0(n898[11])) /* synthesis syn_instantiated=1 */ ;
    IB CE1_pad (.I(CE1), .O(CE1_c));
    LUT4 i23813_3_lut (.A(B_int_adj_661[12]), .B(A_int_adj_660[12]), .C(diffExpAB_adj_668[8]), 
         .Z(efectFracB_adj_666[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23813_3_lut.init = 16'hcaca;
    LUT4 i23789_3_lut (.A(B_int_adj_661[10]), .B(A_int_adj_660[10]), .C(diffExpAB_adj_668[8]), 
         .Z(efectFracB_adj_666[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23789_3_lut.init = 16'hcaca;
    LUT4 i23807_3_lut (.A(B_int_adj_661[11]), .B(A_int_adj_660[11]), .C(diffExpAB_adj_668[8]), 
         .Z(efectFracB_adj_666[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23807_3_lut.init = 16'hcaca;
    \output  output0 (.writeout({writeout}), .new_data(new_data), .SDA_c(SDA_c), 
            .n23639(n23639), .output_new(output_new), .GND_net(inputNumber[31]), 
            .n3988(n3980[0]), .mlp_done(mlp_done), .n28181(n28181), .\mlp_outputs[0] ({\mlp_outputs[0] }), 
            .\mlp_outputs[1] ({\mlp_outputs[1] }), .n66628(n66628), .n73802(n73802));
    LUT4 i23811_3_lut (.A(B_int_adj_661[12]), .B(n480_adj_701[15]), .C(n73825), 
         .Z(frac_adj_677[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23811_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_721_4_lut (.A(B_int_adj_661[10]), .B(n35407), .C(n73825), 
         .D(n70693), .Z(n70691)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_721_4_lut.init = 16'hffca;
    LUT4 i23797_3_lut_rep_722 (.A(B_int_adj_661[10]), .B(n35407), .C(n73825), 
         .Z(n70692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23797_3_lut_rep_722.init = 16'hcaca;
    FD1S1A dlatchrs_7_i1 (.D(writeout[0]), .CK(output_new), .Q(write_data[0]));
    defparam dlatchrs_7_i1.GSR = "DISABLED";
    LUT4 i23796_3_lut (.A(A_int_adj_660[10]), .B(n451_adj_700[13]), .C(n70727), 
         .Z(n35407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23796_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n42939), .B(n42934), .C(n73833), .D(n73837), .Z(FP_Z_int_adj_729[22])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 i24141_3_lut (.A(B_int[3]), .B(A_int[3]), .C(diffExpAB[8]), .Z(n73827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24141_3_lut.init = 16'hcaca;
    LUT4 i6_3_lut (.A(n73827), .B(n70834), .C(diffExp[4]), .Z(n5[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6_3_lut.init = 16'hcaca;
    LUT4 i24011_3_lut (.A(B_int[2]), .B(A_int[2]), .C(diffExpAB[8]), .Z(efectFracB[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24011_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(n42939), .B(exp_final[7]), .Z(n984[7])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i6_3_lut_adj_986 (.A(efectFracB[5]), .B(efectFracB[21]), .C(diffExp[4]), 
         .Z(n5[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6_3_lut_adj_986.init = 16'hcaca;
    LUT4 i23999_3_lut (.A(B_int[4]), .B(A_int[4]), .C(diffExpAB[8]), .Z(efectFracB[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23999_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_987 (.A(n42939), .B(exp_final[6]), .Z(n984[6])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_987.init = 16'h8888;
    LUT4 i24248_3_lut (.A(B_int[9]), .B(A_int[9]), .C(diffExpAB[8]), .Z(efectFracB[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24248_3_lut.init = 16'hcaca;
    LUT4 i24128_3_lut (.A(B_int[10]), .B(A_int[10]), .C(diffExpAB[8]), 
         .Z(efectFracB[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24128_3_lut.init = 16'hcaca;
    LUT4 i24249_3_lut (.A(B_int[11]), .B(A_int[11]), .C(diffExpAB[8]), 
         .Z(efectFracB[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24249_3_lut.init = 16'hcaca;
    LUT4 i24152_3_lut (.A(efectFracB[14]), .B(n70834), .C(n70835), .Z(n19214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24152_3_lut.init = 16'hcaca;
    loadWeight loadWeight0 (.sram_address_A({sram_address_A}), .clock(clock), 
            .n4445(n73830), .sram_input_A({sram_input_A}), .ramDataIn({ramDataIn}), 
            .sram_ready_A(sram_ready_A), .SDA_c(SDA_c), .n73801(n73801), 
            .n1682(n1682), .n1673(n1670[1]), .n73802(n73802), .n39(n39), 
            .n23939(n23939), .GND_net(inputNumber[31]));
    LUT4 i1_2_lut_adj_988 (.A(n42939), .B(exp_final[5]), .Z(n984[5])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_988.init = 16'h8888;
    LUT4 i1_2_lut_adj_989 (.A(n42939), .B(exp_final[4]), .Z(n984[4])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_989.init = 16'h8888;
    LUT4 i1_2_lut_adj_990 (.A(n42939), .B(exp_final[3]), .Z(n984[3])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_990.init = 16'h8888;
    receiver receiver0 (.clock(clock), .SDA_c(SDA_c), .read_data({read_data}), 
            .ramDataIn({ramDataIn}), .count({Open_0, Open_1, Open_2, 
            Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, Open_9, 
            Open_10, Open_11, Open_12, Open_13, Open_14, Open_15, 
            Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, 
            Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, 
            Open_28, Open_29, count[1:0]}), .n63477(n63477), .new_data(new_data), 
            .n25(n73840), .n70855(n70855), .GND_net(inputNumber[31]));
    LUT4 i14337_3_lut (.A(prod[22]), .B(prod[23]), .C(prod[47]), .Z(frac_norm[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14337_3_lut.init = 16'hcaca;
    LUT4 i24235_3_lut (.A(B_int[18]), .B(A_int[18]), .C(diffExpAB[8]), 
         .Z(efectFracB[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24235_3_lut.init = 16'hcaca;
    VLO i1 (.Z(inputNumber[31]));
    PUR PUR_INST (.PUR(inputNumber[2]));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i24246_3_lut (.A(B_int[13]), .B(A_int[13]), .C(diffExpAB[8]), 
         .Z(efectFracB[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24246_3_lut.init = 16'hcaca;
    LUT4 i24000_3_lut (.A(B_int[17]), .B(A_int[17]), .C(diffExpAB[8]), 
         .Z(efectFracB[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24000_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut (.A(prod[23]), .B(prod[24]), .C(prod[47]), .Z(frac_norm[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 i14326_3_lut (.A(prod[25]), .B(prod[26]), .C(prod[47]), .Z(frac_norm[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14326_3_lut.init = 16'hcaca;
    LUT4 i14332_3_lut (.A(prod[24]), .B(prod[25]), .C(prod[47]), .Z(frac_norm[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14332_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_991 (.A(n42939), .B(exp_final[2]), .Z(n984[2])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_991.init = 16'h8888;
    LUT4 i24147_3_lut (.A(B_int[12]), .B(A_int[12]), .C(diffExpAB[8]), 
         .Z(efectFracB[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24147_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_992 (.A(n42939), .B(exp_final[1]), .Z(n984[1])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_992.init = 16'h8888;
    LUT4 i1_2_lut_adj_993 (.A(n42939), .B(exp_final[0]), .Z(n984[0])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_993.init = 16'h8888;
    LUT4 i14336_3_lut (.A(prod[27]), .B(prod[28]), .C(prod[47]), .Z(frac_norm[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14336_3_lut.init = 16'hcaca;
    LUT4 i24016_3_lut (.A(B_int[16]), .B(A_int[16]), .C(diffExpAB[8]), 
         .Z(efectFracB[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24016_3_lut.init = 16'hcaca;
    LUT4 i15_1_lut (.A(prod[47]), .Z(n73831)) /* synthesis lut_function=(!(A)) */ ;
    defparam i15_1_lut.init = 16'h5555;
    spi2 spi0 (.clock(clock), .new_data(new_data), .GND_net(inputNumber[31]), 
         .VCC_net(inputNumber[2]), .CE1_c(CE1_c), .spi_mosi_oe(spi_mosi_oe), 
         .spi_mosi_o(spi_mosi_o), .spi_miso_oe(spi_miso_oe), .spi_miso_o(spi_miso_o), 
         .spi_clk_oe(spi_clk_oe), .spi_clk_o(spi_clk_o), .spi_mosi_i(spi_mosi_i), 
         .spi_miso_i(spi_miso_i), .spi_clk_i(spi_clk_i), .read_data({read_data}), 
         .write_data({write_data}), .n63477(n63477), .n25(n73840), .n39(n39), 
         .\count[0] (count[0]), .\count[1] (count[1]), .n23939(n23939), 
         .n70855(n70855));
    LUT4 i15162_3_lut (.A(prod[28]), .B(prod[29]), .C(prod[47]), .Z(frac_norm[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15162_3_lut.init = 16'hcaca;
    LUT4 i15173_3_lut (.A(prod[31]), .B(prod[32]), .C(prod[47]), .Z(frac_norm[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15173_3_lut.init = 16'hcaca;
    LUT4 i15174_3_lut (.A(prod[30]), .B(prod[31]), .C(prod[47]), .Z(frac_norm[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15174_3_lut.init = 16'hcaca;
    LUT4 i15170_3_lut (.A(prod[33]), .B(prod[34]), .C(prod[47]), .Z(frac_norm[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15170_3_lut.init = 16'hcaca;
    LUT4 i15171_3_lut (.A(prod[32]), .B(prod[33]), .C(prod[47]), .Z(frac_norm[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15171_3_lut.init = 16'hcaca;
    pr pr0 (.n3946(n3942[0]), .clock(clock), .n23661(n23661), .SDA_c(SDA_c), 
       .n73801(n73801), .weight_done(weight_done), .n1682(n1682), .n73802(n73802), 
       .\state[0] (state_adj_642[0]), .n3961(n3961), .n3944(n3942[2]), 
       .n22106(n22106));
    LUT4 i14338_3_lut (.A(prod[35]), .B(prod[36]), .C(prod[47]), .Z(frac_norm[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14338_3_lut.init = 16'hcaca;
    LUT4 i14327_3_lut (.A(prod[34]), .B(prod[35]), .C(prod[47]), .Z(frac_norm[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14327_3_lut.init = 16'hcaca;
    LUT4 i14330_3_lut (.A(prod[36]), .B(prod[37]), .C(prod[47]), .Z(frac_norm[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14330_3_lut.init = 16'hcaca;
    LUT4 i14331_3_lut (.A(prod[40]), .B(prod[41]), .C(prod[47]), .Z(frac_norm[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14331_3_lut.init = 16'hcaca;
    float_alu float_alu0 (.n1151(n1148[5]), .n1156(n1148[0]), .\float_alu_mode[1] (float_alu_mode[1]), 
            .\float_alu_mode[2] (float_alu_mode[2]), .float_alu_c({float_alu_c}), 
            .clock(clock), .n70744(n70744), .n70778(n70778), .SDA_c(SDA_c), 
            .n70716(n70716), .n24013(n24013), .n63113(n63113), .n63130(n63130), 
            .float_alu_b({float_alu_b}), .n62900(n62900), .n124(n73838), 
            .float_alu_ready(float_alu_ready), .n70866(n70866), .n2050(n2022[36]), 
            .n4617(n4617), .n2084(n2022[2]), .n15113(n15113), .n2072(n2022[14]), 
            .n4599(n4599), .n1155(n1148[1]), .n70822(n70822), .n2036(n2022[50]), 
            .n2086(n2022[0]), .n23655(n23655), .n23979(n23979), .n73809(n73809), 
            .n70788(n70788), .n73818(n73818), .n2082(n2022[4]), .n23653(n23653), 
            .n45598(n45598), .n63068(n63068), .n62958(n62958), .n66522(n66522), 
            .n66524(n66524), .n63156(n63156), .n63069(n63069), .n63070(n63070), 
            .n62961(n62961), .n63102(n63102), .n63103(n63103), .n63104(n63104), 
            .n63106(n63106), .n63105(n63105), .n63107(n63107), .n63114(n63114), 
            .n63109(n63109), .n63115(n63115), .n63116(n63116), .n63120(n63120), 
            .n63122(n63122), .n63128(n63128), .n63131(n63131), .n63139(n63139), 
            .n63147(n63147), .n63150(n63150), .n62964(n62964), .n62966(n62966), 
            .n1673(n1670[1]), .n4445(n73830), .n27939(n27939), .n23942(n23942), 
            .n63112(n63112), .n63111(n63111), .n70816(n70816), .GND_net(inputNumber[31]), 
            .n42934(n42934), .n61(n73825), .\A_int[10] (A_int_adj_660[10]), 
            .\B_int[10] (B_int_adj_661[10]), .n70727(n70727), .\A_int[11] (A_int_adj_660[11]), 
            .\B_int[11] (B_int_adj_661[11]), .\A_int[12] (A_int_adj_660[12]), 
            .\B_int[12] (B_int_adj_661[12]), .n70692(n70692), .\frac[15] (frac_adj_677[15]), 
            .n70693(n70693), .\diffExpAB[8] (diffExpAB_adj_668[8]), .n493(n480_adj_701[15]), 
            .n466(n451_adj_700[13]), .n70691(n70691), .\efectFracB[13] (efectFracB_adj_666[13]), 
            .\efectFracB[15] (efectFracB_adj_666[15]), .\efectFracB[14] (efectFracB_adj_666[14]), 
            .\B_int[12]_adj_2 (B_int_adj_725[12]), .\B_int[13] (B_int_adj_725[13]), 
            .\B_int[15] (B_int_adj_725[15]), .\B_int[8] (B_int_adj_725[8]), 
            .\A_int[2] (A_int_adj_724[2]), .\A_int[3] (A_int_adj_724[3]), 
            .\A_int[6] (A_int_adj_724[6]), .\A_int[7] (A_int_adj_724[7]), 
            .\A_int[4] (A_int_adj_724[4]), .\A_int[5] (A_int_adj_724[5]), 
            .\B_int[0] (B_int_adj_725[0]), .\A_int[0] (A_int_adj_724[0]), 
            .\A_int[11]_adj_3 (A_int_adj_724[11]), .\A_int[12]_adj_4 (A_int_adj_724[12]), 
            .\A_int[13] (A_int_adj_724[13]), .\A_int[15] (A_int_adj_724[15]), 
            .\A_int[17] (A_int_adj_724[17]), .\A_int[16] (A_int_adj_724[16]), 
            .\A_int[18] (A_int_adj_724[18]), .\A_int[19] (A_int_adj_724[19]), 
            .\A_int[14] (A_int_adj_724[14]), .n4(n73833), .n41520(n41520), 
            .\A_int[1] (A_int_adj_724[1]), .\A_int[10]_adj_5 (A_int_adj_724[10]), 
            .\A_int[9] (A_int_adj_724[9]), .\A_int[22] (A_int_adj_724[22]), 
            .\A_int[21] (A_int_adj_724[21]), .\A_int[8] (A_int_adj_724[8]), 
            .\A_int[20] (A_int_adj_724[20]), .n22310(n22310), .\B_int[11]_adj_6 (B_int_adj_725[11]), 
            .\B_int[14] (B_int_adj_725[14]), .\B_int[10]_adj_7 (B_int_adj_725[10]), 
            .\B_int[9] (B_int_adj_725[9]), .\B_int[19] (B_int_adj_725[19]), 
            .\B_int[18] (B_int_adj_725[18]), .\B_int[20] (B_int_adj_725[20]), 
            .\B_int[21] (B_int_adj_725[21]), .\B_int[7] (B_int_adj_725[7]), 
            .n22437(n22437), .\prod[47] (prod[47]), .n66955(n66955), .n67025(n67025), 
            .n67007(n67007), .\prod[45] (prod[45]), .\prod[46] (prod[46]), 
            .\prod[28] (prod[28]), .\prod[33] (prod[33]), .\prod[40] (prod[40]), 
            .\prod[22] (prod[22]), .\prod[24] (prod[24]), .\prod[25] (prod[25]), 
            .\prod[23] (prod[23]), .\prod[26] (prod[26]), .\prod[41] (prod[41]), 
            .\prod[34] (prod[34]), .\prod[37] (prod[37]), .\prod[27] (prod[27]), 
            .\prod[39] (prod[39]), .\prod[29] (prod[29]), .\prod[35] (prod[35]), 
            .\prod[36] (prod[36]), .\prod[31] (prod[31]), .\prod[32] (prod[32]), 
            .\prod[43] (prod[43]), .\prod[30] (prod[30]), .\prod[38] (prod[38]), 
            .\prod[42] (prod[42]), .\prod[44] (prod[44]), .n42939(n42939), 
            .n25571(n25571), .\frac_norm[20] (frac_norm[20]), .\frac_norm[16] (frac_norm[16]), 
            .\frac_norm[14] (frac_norm[14]), .\frac_norm[15] (frac_norm[15]), 
            .\frac_norm[12] (frac_norm[12]), .\frac_norm[13] (frac_norm[13]), 
            .\frac_norm[10] (frac_norm[10]), .\frac_norm[11] (frac_norm[11]), 
            .\frac_norm[8] (frac_norm[8]), .n15(n73831), .\B_int[17] (B_int_adj_725[17]), 
            .\B_int[16] (B_int_adj_725[16]), .\B_int[22] (B_int_adj_725[22]), 
            .\frac_norm[7] (frac_norm[7]), .n984({n984}), .\B_int[3] (B_int_adj_725[3]), 
            .\B_int[1] (B_int_adj_725[1]), .\B_int[2] (B_int_adj_725[2]), 
            .\frac_norm[4] (frac_norm[4]), .\frac_norm[5] (frac_norm[5]), 
            .\frac_norm[3] (frac_norm[3]), .\frac_norm[2] (frac_norm[2]), 
            .exp_final({exp_final}), .\FP_Z_int[22] (FP_Z_int_adj_729[22]), 
            .\B_int[6] (B_int_adj_725[6]), .\B_int[5] (B_int_adj_725[5]), 
            .\B_int[4] (B_int_adj_725[4]), .n6(n73837), .\prod[21] (prod[21]), 
            .VCC_net(inputNumber[2]), .\buf_x[89] (buf_x_adj_1109[89]), 
            .\buf_x[87] (buf_x_adj_1109[87]), .\buf_x[88] (buf_x_adj_1109[88]), 
            .\buf_x[85] (buf_x_adj_1109[85]), .\buf_x[86] (buf_x_adj_1109[86]), 
            .\buf_x[83] (buf_x_adj_1109[83]), .\buf_x[84] (buf_x_adj_1109[84]), 
            .\buf_r[89] (buf_r_adj_1110[89]), .\buf_r[87] (buf_r_adj_1110[87]), 
            .\buf_r[88] (buf_r_adj_1110[88]), .\buf_r[85] (buf_r_adj_1110[85]), 
            .\buf_r[86] (buf_r_adj_1110[86]), .\buf_r[83] (buf_r_adj_1110[83]), 
            .\buf_r[84] (buf_r_adj_1110[84]), .\A_int[11]_adj_8 (A_int[11]), 
            .\B_int[11]_adj_9 (B_int[11]), .\A_int[10]_adj_10 (A_int[10]), 
            .\B_int[10]_adj_11 (B_int[10]), .\A_int[13]_adj_12 (A_int[13]), 
            .\B_int[13]_adj_13 (B_int[13]), .\A_int[12]_adj_14 (A_int[12]), 
            .\B_int[12]_adj_15 (B_int[12]), .\A_int[17]_adj_16 (A_int[17]), 
            .\B_int[17]_adj_17 (B_int[17]), .\A_int[16]_adj_18 (A_int[16]), 
            .\B_int[16]_adj_19 (B_int[16]), .\A_int[18]_adj_20 (A_int[18]), 
            .\B_int[18]_adj_21 (B_int[18]), .\A_int[2]_adj_22 (A_int[2]), 
            .\B_int[2]_adj_23 (B_int[2]), .\B_int[3]_adj_24 (B_int[3]), 
            .\A_int[9]_adj_25 (A_int[9]), .\A_int[7]_adj_26 (A_int[7]), 
            .\A_int[4]_adj_27 (A_int[4]), .\A_int[3]_adj_28 (A_int[3]), 
            .\B_int[9]_adj_29 (B_int[9]), .\B_int[7]_adj_30 (B_int[7]), 
            .\B_int[4]_adj_31 (B_int[4]), .\diffExpAB[8]_adj_32 (diffExpAB[8]), 
            .\diffExp[4] (diffExp[4]), .n70835(n70835), .n70834(n70834), 
            .n70833(n70833), .\efectFracB[21] (efectFracB[21]), .\efectFracB[20] (efectFracB[20]), 
            .\efectFracB[19] (efectFracB[19]), .\efectFracB[15]_adj_33 (efectFracB[15]), 
            .\efectFracB[16] (efectFracB[16]), .n19214(n19214), .n28(n5[5]), 
            .n70771(n70771), .n9(n73827), .\efectFracB[14]_adj_34 (efectFracB[14]), 
            .\efectFracB[7] (efectFracB[7]), .\efectFracB[5] (efectFracB[5]), 
            .\efectFracB[12] (efectFracB[12]), .n70820(n70820), .\efectFracB[13]_adj_35 (efectFracB[13]), 
            .n27(n5[6]), .n70740(n70740), .n55(n37_adj_763[10]));
    LUT4 m1_lut (.Z(n73802)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    test test0 (.sram_address_B({sram_address_B}), .clock(clock), .GND_net(inputNumber[31]), 
         .sram_output_B({sram_output_B}), .n4599(n4599), .float_alu_c({float_alu_c}), 
         .i({Open_30, Open_31, Open_32, Open_33, Open_34, Open_35, 
         Open_36, Open_37, Open_38, Open_39, Open_40, Open_41, Open_42, 
         Open_43, Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, 
         Open_50, i[10], Open_51, Open_52, Open_53, Open_54, Open_55, 
         Open_56, Open_57, i[2:0]}), .n15113(n15113), .n4617(n4617), 
         .n14054(n14053[1]), .n70822(n70822), .\mlp_outputs[0] ({\mlp_outputs[0] }), 
         .\mlp_outputs[1] ({\mlp_outputs[1] }), .n23653(n23653), .SDA_c(SDA_c), 
         .sram_ready_B(sram_ready_B), .n23655(n23655), .weight_done(weight_done), 
         .n2086(n2022[0]), .n70866(n70866), .float_alu_ready(float_alu_ready), 
         .float_alu_b({float_alu_b}), .n927(n898[5]), .n926(n898[6]), 
         .n70778(n70778), .n70788(n70788), .n14050(n14049[1]), .n2889({n2889}), 
         .n3044({n3044}), .n236({n236}), .n61382(n61382), .n63111(n63111), 
         .n23661(n23661), .\float_alu_mode[1] (float_alu_mode[1]), .n27939(n27939), 
         .n63112(n63112), .\i[8] (i[8]), .\i[9] (i[9]), .n929(n898[3]), 
         .n928(n898[4]), .\buf_r[83] (buf_r_adj_1110[83]), .\buf_x[83] (buf_x_adj_1109[83]), 
         .n2082(n2022[4]), .n73818(n73818), .n923(n898[9]), .n922(n898[10]), 
         .\state[0] (state_adj_642[0]), .\float_alu_mode[2] (float_alu_mode[2]), 
         .n1155(n1148[1]), .n124(n73838), .n2036(n2022[50]), .n70816(n70816), 
         .n2050(n2022[36]), .n2072(n2022[14]), .n2084(n2022[2]), .\i[12] (i[12]), 
         .\i[11] (i[11]), .\i[7] (i[7]), .\i[6] (i[6]), .\i[5] (i[5]), 
         .\i[4] (i[4]), .\i[3] (i[3]), .n70716(n70716), .n24013(n24013), 
         .n62900(n62900), .n932(n898[0]), .n930(n898[2]), .n63130(n63130), 
         .\buf_r[84] (buf_r_adj_1110[84]), .\buf_x[84] (buf_x_adj_1109[84]), 
         .\buf_r[85] (buf_r_adj_1110[85]), .\buf_x[85] (buf_x_adj_1109[85]), 
         .\buf_r[86] (buf_r_adj_1110[86]), .\buf_x[86] (buf_x_adj_1109[86]), 
         .\buf_r[87] (buf_r_adj_1110[87]), .\buf_x[87] (buf_x_adj_1109[87]), 
         .\buf_r[88] (buf_r_adj_1110[88]), .\buf_x[88] (buf_x_adj_1109[88]), 
         .\buf_r[89] (buf_r_adj_1110[89]), .\buf_x[89] (buf_x_adj_1109[89]), 
         .n63113(n63113), .mlp_done(mlp_done), .n73801(n73801), .n3946(n3942[0]), 
         .n3944(n3942[2]), .n22106(n22106), .n3961(n3961), .n62966(n62966), 
         .n62964(n62964), .n63150(n63150), .n63147(n63147), .n63139(n63139), 
         .n63131(n63131), .n63128(n63128), .n63122(n63122), .n63120(n63120), 
         .n63116(n63116), .n63115(n63115), .n63109(n63109), .n63114(n63114), 
         .n63107(n63107), .n63105(n63105), .n63106(n63106), .n63104(n63104), 
         .n63103(n63103), .n63102(n63102), .n62961(n62961), .n63070(n63070), 
         .n63069(n63069), .n63156(n63156), .n66524(n66524), .n66522(n66522), 
         .n62958(n62958), .n63068(n63068), .n70867(n70867), .n921(n898[11]), 
         .n23942(n23942), .n3988(n3980[0]), .n28181(n28181), .n66628(n66628), 
         .n23639(n23639), .n1156(n1148[0]), .n73809(n73809), .n45598(n45598), 
         .n931(n898[1]), .n925(n898[7]), .n924(n898[8]));
    LUT4 i49744_1_lut (.A(n236[0]), .Z(n61382)) /* synthesis lut_function=(!(A)) */ ;
    defparam i49744_1_lut.init = 16'h5555;
    sram_dp sram_dp0 (.sram_input_A({sram_input_A}), .GND_net(inputNumber[31]), 
            .sram_address_A({sram_address_A}), .sram_address_B({sram_address_B}), 
            .clock(clock), .sram_ready_A(sram_ready_A), .sram_ready_B(sram_ready_B), 
            .VCC_net(inputNumber[2]), .SDA_c(SDA_c), .sram_output_B({sram_output_B}));
    
endmodule
//
// Verilog Description of module \output 
//

module \output  (writeout, new_data, SDA_c, n23639, output_new, GND_net, 
            n3988, mlp_done, n28181, \mlp_outputs[0] , \mlp_outputs[1] , 
            n66628, n73802);
    output [7:0]writeout;
    input new_data;
    input SDA_c;
    input n23639;
    output output_new;
    input GND_net;
    output n3988;
    input mlp_done;
    output n28181;
    input [31:0]\mlp_outputs[0] ;
    input [31:0]\mlp_outputs[1] ;
    input n66628;
    input n73802;
    
    wire [31:0]dat_reg;   // c:/users/yisong/documents/new/mlp/output.vhd(29[8:15])
    wire [31:0]k;   // c:/users/yisong/documents/new/mlp/output.vhd(28[8:9])
    wire n73802 /* synthesis nomerge= */ ;
    
    wire n23638;
    wire [7:0]n13501;
    wire [31:0]n8;
    
    wire n23657;
    wire [7:0]n3980;
    
    wire n62629;
    wire [31:0]n134;
    
    wire n62628, n62627, n62626, n62625, n62624, n62623, n62622, 
        n62621, n62620, n62619, n62618, n62617, n62616, n62615, 
        n38, n52, n48, n55, n42, n54, n60, n41, n50, n58, 
        n62, n49, n28182;
    wire [7:0]n13471;
    wire [7:0]n13481;
    
    wire n13490;
    
    FD1P3DX DataOut_i0_i0 (.D(n13501[0]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[0]));
    defparam DataOut_i0_i0.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i0 (.D(n8[0]), .SP(n23639), .CK(new_data), .Q(dat_reg[0]));
    defparam dat_reg_i0_i0.GSR = "DISABLED";
    FD1P3DX output_new_34 (.D(n3980[1]), .SP(n23657), .CK(new_data), .CD(SDA_c), 
            .Q(output_new));
    defparam output_new_34.GSR = "DISABLED";
    CCU2D k_4662_add_4_32 (.A0(k[30]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62629), 
          .S0(n134[30]), .S1(n134[31]));
    defparam k_4662_add_4_32.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_32.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_32.INJECT1_0 = "NO";
    defparam k_4662_add_4_32.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_30 (.A0(k[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62628), 
          .COUT(n62629), .S0(n134[28]), .S1(n134[29]));
    defparam k_4662_add_4_30.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_30.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_30.INJECT1_0 = "NO";
    defparam k_4662_add_4_30.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_28 (.A0(k[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62627), 
          .COUT(n62628), .S0(n134[26]), .S1(n134[27]));
    defparam k_4662_add_4_28.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_28.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_28.INJECT1_0 = "NO";
    defparam k_4662_add_4_28.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_26 (.A0(k[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62626), 
          .COUT(n62627), .S0(n134[24]), .S1(n134[25]));
    defparam k_4662_add_4_26.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_26.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_26.INJECT1_0 = "NO";
    defparam k_4662_add_4_26.INJECT1_1 = "NO";
    FD1P3BX state_FSM__i1 (.D(n3980[4]), .SP(mlp_done), .CK(new_data), 
            .PD(SDA_c), .Q(n3988));
    defparam state_FSM__i1.GSR = "DISABLED";
    CCU2D k_4662_add_4_24 (.A0(k[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62625), 
          .COUT(n62626), .S0(n134[22]), .S1(n134[23]));
    defparam k_4662_add_4_24.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_24.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_24.INJECT1_0 = "NO";
    defparam k_4662_add_4_24.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_22 (.A0(k[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62624), 
          .COUT(n62625), .S0(n134[20]), .S1(n134[21]));
    defparam k_4662_add_4_22.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_22.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_22.INJECT1_0 = "NO";
    defparam k_4662_add_4_22.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_20 (.A0(k[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62623), 
          .COUT(n62624), .S0(n134[18]), .S1(n134[19]));
    defparam k_4662_add_4_20.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_20.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_20.INJECT1_0 = "NO";
    defparam k_4662_add_4_20.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_18 (.A0(k[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62622), 
          .COUT(n62623), .S0(n134[16]), .S1(n134[17]));
    defparam k_4662_add_4_18.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_18.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_18.INJECT1_0 = "NO";
    defparam k_4662_add_4_18.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_16 (.A0(k[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62621), 
          .COUT(n62622), .S0(n134[14]), .S1(n134[15]));
    defparam k_4662_add_4_16.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_16.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_16.INJECT1_0 = "NO";
    defparam k_4662_add_4_16.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_14 (.A0(k[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62620), 
          .COUT(n62621), .S0(n134[12]), .S1(n134[13]));
    defparam k_4662_add_4_14.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_14.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_14.INJECT1_0 = "NO";
    defparam k_4662_add_4_14.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_12 (.A0(k[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62619), 
          .COUT(n62620), .S0(n134[10]), .S1(n134[11]));
    defparam k_4662_add_4_12.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_12.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_12.INJECT1_0 = "NO";
    defparam k_4662_add_4_12.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_10 (.A0(k[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62618), 
          .COUT(n62619), .S0(n134[8]), .S1(n134[9]));
    defparam k_4662_add_4_10.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_10.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_10.INJECT1_0 = "NO";
    defparam k_4662_add_4_10.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_8 (.A0(k[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62617), 
          .COUT(n62618), .S0(n134[6]), .S1(n134[7]));
    defparam k_4662_add_4_8.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_8.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_8.INJECT1_0 = "NO";
    defparam k_4662_add_4_8.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_6 (.A0(k[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62616), 
          .COUT(n62617), .S0(n134[4]), .S1(n134[5]));
    defparam k_4662_add_4_6.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_6.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_6.INJECT1_0 = "NO";
    defparam k_4662_add_4_6.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_4 (.A0(k[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(k[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62615), 
          .COUT(n62616), .S0(n134[2]), .S1(n134[3]));
    defparam k_4662_add_4_4.INIT0 = 16'hfaaa;
    defparam k_4662_add_4_4.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_4.INJECT1_0 = "NO";
    defparam k_4662_add_4_4.INJECT1_1 = "NO";
    CCU2D k_4662_add_4_2 (.A0(n3980[4]), .B0(k[0]), .C0(GND_net), .D0(GND_net), 
          .A1(k[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62615), 
          .S1(n134[1]));
    defparam k_4662_add_4_2.INIT0 = 16'h7000;
    defparam k_4662_add_4_2.INIT1 = 16'hfaaa;
    defparam k_4662_add_4_2.INJECT1_0 = "NO";
    defparam k_4662_add_4_2.INJECT1_1 = "NO";
    FD1P3DX DataOut_i0_i7 (.D(n13501[7]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[7]));
    defparam DataOut_i0_i7.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i6 (.D(n13501[6]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[6]));
    defparam DataOut_i0_i6.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i5 (.D(n13501[5]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[5]));
    defparam DataOut_i0_i5.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i4 (.D(n13501[4]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[4]));
    defparam DataOut_i0_i4.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i3 (.D(n13501[3]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[3]));
    defparam DataOut_i0_i3.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i2 (.D(n13501[2]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[2]));
    defparam DataOut_i0_i2.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i1 (.D(n13501[1]), .SP(n23638), .CK(new_data), 
            .CD(SDA_c), .Q(writeout[1]));
    defparam DataOut_i0_i1.GSR = "DISABLED";
    LUT4 i6_2_lut (.A(k[14]), .B(k[25]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(k[10]), .B(k[0]), .C(k[21]), .D(k[23]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i16_2_lut (.A(k[3]), .B(k[20]), .Z(n48)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i16_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(k[5]), .B(k[7]), .C(k[6]), .D(k[24]), .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(k[29]), .B(k[11]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(k[19]), .B(k[8]), .C(k[2]), .D(k[16]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i28_4_lut (.A(n55), .B(k[1]), .C(n48), .D(k[4]), .Z(n60)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i28_4_lut.init = 16'hfffb;
    LUT4 i9_2_lut (.A(k[9]), .B(k[26]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(n3988), .B(mlp_done), .C(n3980[1]), .Z(n23657)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut.init = 16'hc8c8;
    LUT4 i18_4_lut (.A(k[12]), .B(k[27]), .C(k[17]), .D(k[28]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(k[22]), .B(n52), .C(n38), .D(k[30]), .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(k[18]), .B(k[13]), .C(k[31]), .D(k[15]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i31_4_lut (.A(n49), .B(n62), .C(n58), .D(n50), .Z(n28181)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 mux_7_Mux_0_i1_3_lut (.A(\mlp_outputs[0] [0]), .B(\mlp_outputs[1] [0]), 
         .C(k[0]), .Z(n8[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_0_i1_3_lut.init = 16'hcaca;
    FD1P3DX k_4662__i0 (.D(n134[0]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[0]));
    defparam k_4662__i0.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i31 (.D(n8[31]), .SP(n23639), .CK(new_data), .Q(dat_reg[31]));
    defparam dat_reg_i0_i31.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i30 (.D(n8[30]), .SP(n23639), .CK(new_data), .Q(dat_reg[30]));
    defparam dat_reg_i0_i30.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i29 (.D(n8[29]), .SP(n23639), .CK(new_data), .Q(dat_reg[29]));
    defparam dat_reg_i0_i29.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i28 (.D(n8[28]), .SP(n23639), .CK(new_data), .Q(dat_reg[28]));
    defparam dat_reg_i0_i28.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i27 (.D(n8[27]), .SP(n23639), .CK(new_data), .Q(dat_reg[27]));
    defparam dat_reg_i0_i27.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i26 (.D(n8[26]), .SP(n23639), .CK(new_data), .Q(dat_reg[26]));
    defparam dat_reg_i0_i26.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i25 (.D(n8[25]), .SP(n23639), .CK(new_data), .Q(dat_reg[25]));
    defparam dat_reg_i0_i25.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i24 (.D(n8[24]), .SP(n23639), .CK(new_data), .Q(dat_reg[24]));
    defparam dat_reg_i0_i24.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i23 (.D(n8[23]), .SP(n23639), .CK(new_data), .Q(dat_reg[23]));
    defparam dat_reg_i0_i23.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i22 (.D(n8[22]), .SP(n23639), .CK(new_data), .Q(dat_reg[22]));
    defparam dat_reg_i0_i22.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i21 (.D(n8[21]), .SP(n23639), .CK(new_data), .Q(dat_reg[21]));
    defparam dat_reg_i0_i21.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i20 (.D(n8[20]), .SP(n23639), .CK(new_data), .Q(dat_reg[20]));
    defparam dat_reg_i0_i20.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i19 (.D(n8[19]), .SP(n23639), .CK(new_data), .Q(dat_reg[19]));
    defparam dat_reg_i0_i19.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i18 (.D(n8[18]), .SP(n23639), .CK(new_data), .Q(dat_reg[18]));
    defparam dat_reg_i0_i18.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i17 (.D(n8[17]), .SP(n23639), .CK(new_data), .Q(dat_reg[17]));
    defparam dat_reg_i0_i17.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i16 (.D(n8[16]), .SP(n23639), .CK(new_data), .Q(dat_reg[16]));
    defparam dat_reg_i0_i16.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i15 (.D(n8[15]), .SP(n23639), .CK(new_data), .Q(dat_reg[15]));
    defparam dat_reg_i0_i15.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i14 (.D(n8[14]), .SP(n23639), .CK(new_data), .Q(dat_reg[14]));
    defparam dat_reg_i0_i14.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i13 (.D(n8[13]), .SP(n23639), .CK(new_data), .Q(dat_reg[13]));
    defparam dat_reg_i0_i13.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i12 (.D(n8[12]), .SP(n23639), .CK(new_data), .Q(dat_reg[12]));
    defparam dat_reg_i0_i12.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i11 (.D(n8[11]), .SP(n23639), .CK(new_data), .Q(dat_reg[11]));
    defparam dat_reg_i0_i11.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i10 (.D(n8[10]), .SP(n23639), .CK(new_data), .Q(dat_reg[10]));
    defparam dat_reg_i0_i10.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i9 (.D(n8[9]), .SP(n23639), .CK(new_data), .Q(dat_reg[9]));
    defparam dat_reg_i0_i9.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i8 (.D(n8[8]), .SP(n23639), .CK(new_data), .Q(dat_reg[8]));
    defparam dat_reg_i0_i8.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i7 (.D(n8[7]), .SP(n23639), .CK(new_data), .Q(dat_reg[7]));
    defparam dat_reg_i0_i7.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i6 (.D(n8[6]), .SP(n23639), .CK(new_data), .Q(dat_reg[6]));
    defparam dat_reg_i0_i6.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i5 (.D(n8[5]), .SP(n23639), .CK(new_data), .Q(dat_reg[5]));
    defparam dat_reg_i0_i5.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i4 (.D(n8[4]), .SP(n23639), .CK(new_data), .Q(dat_reg[4]));
    defparam dat_reg_i0_i4.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i3 (.D(n8[3]), .SP(n23639), .CK(new_data), .Q(dat_reg[3]));
    defparam dat_reg_i0_i3.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i2 (.D(n8[2]), .SP(n23639), .CK(new_data), .Q(dat_reg[2]));
    defparam dat_reg_i0_i2.GSR = "DISABLED";
    FD1P3AX dat_reg_i0_i1 (.D(n8[1]), .SP(n23639), .CK(new_data), .Q(dat_reg[1]));
    defparam dat_reg_i0_i1.GSR = "DISABLED";
    LUT4 i1_3_lut_adj_982 (.A(mlp_done), .B(n3988), .C(n3980[5]), .Z(n23638)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_982.init = 16'h0202;
    LUT4 i1_2_lut (.A(n3988), .B(n28181), .Z(n28182)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    FD1P3DX state_FSM__i2 (.D(n28182), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(n3980[1]));
    defparam state_FSM__i2.GSR = "DISABLED";
    FD1P3DX state_FSM__i3 (.D(n3980[1]), .SP(mlp_done), .CK(new_data), 
            .CD(SDA_c), .Q(n3980[2]));
    defparam state_FSM__i3.GSR = "DISABLED";
    FD1P3DX state_FSM__i4 (.D(n3980[2]), .SP(mlp_done), .CK(new_data), 
            .CD(SDA_c), .Q(n3980[3]));
    defparam state_FSM__i4.GSR = "DISABLED";
    FD1P3DX state_FSM__i5 (.D(n3980[3]), .SP(mlp_done), .CK(new_data), 
            .CD(SDA_c), .Q(n3980[4]));
    defparam state_FSM__i5.GSR = "DISABLED";
    FD1P3DX state_FSM__i6 (.D(n73802), .SP(n66628), .CK(new_data), .CD(SDA_c), 
            .Q(n3980[5]));
    defparam state_FSM__i6.GSR = "DISABLED";
    FD1P3DX k_4662__i1 (.D(n134[1]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[1]));
    defparam k_4662__i1.GSR = "DISABLED";
    FD1P3DX k_4662__i2 (.D(n134[2]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[2]));
    defparam k_4662__i2.GSR = "DISABLED";
    FD1P3DX k_4662__i3 (.D(n134[3]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[3]));
    defparam k_4662__i3.GSR = "DISABLED";
    FD1P3DX k_4662__i4 (.D(n134[4]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[4]));
    defparam k_4662__i4.GSR = "DISABLED";
    FD1P3DX k_4662__i5 (.D(n134[5]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[5]));
    defparam k_4662__i5.GSR = "DISABLED";
    FD1P3DX k_4662__i6 (.D(n134[6]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[6]));
    defparam k_4662__i6.GSR = "DISABLED";
    FD1P3DX k_4662__i7 (.D(n134[7]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[7]));
    defparam k_4662__i7.GSR = "DISABLED";
    FD1P3DX k_4662__i8 (.D(n134[8]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[8]));
    defparam k_4662__i8.GSR = "DISABLED";
    FD1P3DX k_4662__i9 (.D(n134[9]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[9]));
    defparam k_4662__i9.GSR = "DISABLED";
    FD1P3DX k_4662__i10 (.D(n134[10]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[10]));
    defparam k_4662__i10.GSR = "DISABLED";
    FD1P3DX k_4662__i11 (.D(n134[11]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[11]));
    defparam k_4662__i11.GSR = "DISABLED";
    FD1P3DX k_4662__i12 (.D(n134[12]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[12]));
    defparam k_4662__i12.GSR = "DISABLED";
    FD1P3DX k_4662__i13 (.D(n134[13]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[13]));
    defparam k_4662__i13.GSR = "DISABLED";
    FD1P3DX k_4662__i14 (.D(n134[14]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[14]));
    defparam k_4662__i14.GSR = "DISABLED";
    FD1P3DX k_4662__i15 (.D(n134[15]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[15]));
    defparam k_4662__i15.GSR = "DISABLED";
    FD1P3DX k_4662__i16 (.D(n134[16]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[16]));
    defparam k_4662__i16.GSR = "DISABLED";
    FD1P3DX k_4662__i17 (.D(n134[17]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[17]));
    defparam k_4662__i17.GSR = "DISABLED";
    FD1P3DX k_4662__i18 (.D(n134[18]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[18]));
    defparam k_4662__i18.GSR = "DISABLED";
    FD1P3DX k_4662__i19 (.D(n134[19]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[19]));
    defparam k_4662__i19.GSR = "DISABLED";
    FD1P3DX k_4662__i20 (.D(n134[20]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[20]));
    defparam k_4662__i20.GSR = "DISABLED";
    FD1P3DX k_4662__i21 (.D(n134[21]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[21]));
    defparam k_4662__i21.GSR = "DISABLED";
    FD1P3DX k_4662__i22 (.D(n134[22]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[22]));
    defparam k_4662__i22.GSR = "DISABLED";
    FD1P3DX k_4662__i23 (.D(n134[23]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[23]));
    defparam k_4662__i23.GSR = "DISABLED";
    FD1P3DX k_4662__i24 (.D(n134[24]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[24]));
    defparam k_4662__i24.GSR = "DISABLED";
    FD1P3DX k_4662__i25 (.D(n134[25]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[25]));
    defparam k_4662__i25.GSR = "DISABLED";
    FD1P3DX k_4662__i26 (.D(n134[26]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[26]));
    defparam k_4662__i26.GSR = "DISABLED";
    FD1P3DX k_4662__i27 (.D(n134[27]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[27]));
    defparam k_4662__i27.GSR = "DISABLED";
    FD1P3DX k_4662__i28 (.D(n134[28]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[28]));
    defparam k_4662__i28.GSR = "DISABLED";
    FD1P3DX k_4662__i29 (.D(n134[29]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[29]));
    defparam k_4662__i29.GSR = "DISABLED";
    FD1P3DX k_4662__i30 (.D(n134[30]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[30]));
    defparam k_4662__i30.GSR = "DISABLED";
    FD1P3DX k_4662__i31 (.D(n134[31]), .SP(mlp_done), .CK(new_data), .CD(SDA_c), 
            .Q(k[31]));
    defparam k_4662__i31.GSR = "DISABLED";
    LUT4 mux_7_Mux_1_i1_3_lut (.A(\mlp_outputs[0] [1]), .B(\mlp_outputs[1] [1]), 
         .C(k[0]), .Z(n8[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_1_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_2_i1_3_lut (.A(\mlp_outputs[0] [2]), .B(\mlp_outputs[1] [2]), 
         .C(k[0]), .Z(n8[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_3_i1_3_lut (.A(\mlp_outputs[0] [3]), .B(\mlp_outputs[1] [3]), 
         .C(k[0]), .Z(n8[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_4_i1_3_lut (.A(\mlp_outputs[0] [4]), .B(\mlp_outputs[1] [4]), 
         .C(k[0]), .Z(n8[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_5_i1_3_lut (.A(\mlp_outputs[0] [5]), .B(\mlp_outputs[1] [5]), 
         .C(k[0]), .Z(n8[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_6_i1_3_lut (.A(\mlp_outputs[0] [6]), .B(\mlp_outputs[1] [6]), 
         .C(k[0]), .Z(n8[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_7_i1_3_lut (.A(\mlp_outputs[0] [7]), .B(\mlp_outputs[1] [7]), 
         .C(k[0]), .Z(n8[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_8_i1_3_lut (.A(\mlp_outputs[0] [8]), .B(\mlp_outputs[1] [8]), 
         .C(k[0]), .Z(n8[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_8_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_9_i1_3_lut (.A(\mlp_outputs[0] [9]), .B(\mlp_outputs[1] [9]), 
         .C(k[0]), .Z(n8[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_9_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_10_i1_3_lut (.A(\mlp_outputs[0] [10]), .B(\mlp_outputs[1] [10]), 
         .C(k[0]), .Z(n8[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_10_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_11_i1_3_lut (.A(\mlp_outputs[0] [11]), .B(\mlp_outputs[1] [11]), 
         .C(k[0]), .Z(n8[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_11_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_12_i1_3_lut (.A(\mlp_outputs[0] [12]), .B(\mlp_outputs[1] [12]), 
         .C(k[0]), .Z(n8[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_12_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_13_i1_3_lut (.A(\mlp_outputs[0] [13]), .B(\mlp_outputs[1] [13]), 
         .C(k[0]), .Z(n8[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_13_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_14_i1_3_lut (.A(\mlp_outputs[0] [14]), .B(\mlp_outputs[1] [14]), 
         .C(k[0]), .Z(n8[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_14_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_15_i1_3_lut (.A(\mlp_outputs[0] [15]), .B(\mlp_outputs[1] [15]), 
         .C(k[0]), .Z(n8[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_15_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_16_i1_3_lut (.A(\mlp_outputs[0] [16]), .B(\mlp_outputs[1] [16]), 
         .C(k[0]), .Z(n8[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_16_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_17_i1_3_lut (.A(\mlp_outputs[0] [17]), .B(\mlp_outputs[1] [17]), 
         .C(k[0]), .Z(n8[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_17_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_18_i1_3_lut (.A(\mlp_outputs[0] [18]), .B(\mlp_outputs[1] [18]), 
         .C(k[0]), .Z(n8[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_18_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_19_i1_3_lut (.A(\mlp_outputs[0] [19]), .B(\mlp_outputs[1] [19]), 
         .C(k[0]), .Z(n8[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_19_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_20_i1_3_lut (.A(\mlp_outputs[0] [20]), .B(\mlp_outputs[1] [20]), 
         .C(k[0]), .Z(n8[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_20_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_21_i1_3_lut (.A(\mlp_outputs[0] [21]), .B(\mlp_outputs[1] [21]), 
         .C(k[0]), .Z(n8[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_21_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_22_i1_3_lut (.A(\mlp_outputs[0] [22]), .B(\mlp_outputs[1] [22]), 
         .C(k[0]), .Z(n8[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_22_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_23_i1_3_lut (.A(\mlp_outputs[0] [23]), .B(\mlp_outputs[1] [23]), 
         .C(k[0]), .Z(n8[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_23_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_24_i1_3_lut (.A(\mlp_outputs[0] [24]), .B(\mlp_outputs[1] [24]), 
         .C(k[0]), .Z(n8[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_24_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_25_i1_3_lut (.A(\mlp_outputs[0] [25]), .B(\mlp_outputs[1] [25]), 
         .C(k[0]), .Z(n8[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_25_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_26_i1_3_lut (.A(\mlp_outputs[0] [26]), .B(\mlp_outputs[1] [26]), 
         .C(k[0]), .Z(n8[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_26_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_27_i1_3_lut (.A(\mlp_outputs[0] [27]), .B(\mlp_outputs[1] [27]), 
         .C(k[0]), .Z(n8[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_27_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_28_i1_3_lut (.A(\mlp_outputs[0] [28]), .B(\mlp_outputs[1] [28]), 
         .C(k[0]), .Z(n8[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_28_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_29_i1_3_lut (.A(\mlp_outputs[0] [29]), .B(\mlp_outputs[1] [29]), 
         .C(k[0]), .Z(n8[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_29_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_30_i1_3_lut (.A(\mlp_outputs[0] [30]), .B(\mlp_outputs[1] [30]), 
         .C(k[0]), .Z(n8[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_30_i1_3_lut.init = 16'hcaca;
    LUT4 mux_7_Mux_31_i1_3_lut (.A(\mlp_outputs[0] [31]), .B(\mlp_outputs[1] [31]), 
         .C(k[0]), .Z(n8[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_7_Mux_31_i1_3_lut.init = 16'hcaca;
    LUT4 i49861_2_lut (.A(n3980[4]), .B(k[0]), .Z(n134[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49861_2_lut.init = 16'h6666;
    PFUMX mux_4250_i8 (.BLUT(n13471[7]), .ALUT(n13481[7]), .C0(n13490), 
          .Z(n13501[7]));
    PFUMX mux_4250_i7 (.BLUT(n13471[6]), .ALUT(n13481[6]), .C0(n13490), 
          .Z(n13501[6]));
    LUT4 mux_4246_i1_3_lut (.A(dat_reg[8]), .B(dat_reg[0]), .C(n3980[4]), 
         .Z(n13481[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i1_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i1_3_lut (.A(dat_reg[24]), .B(dat_reg[16]), .C(n3980[2]), 
         .Z(n13471[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i1_3_lut.init = 16'hcaca;
    PFUMX mux_4250_i6 (.BLUT(n13471[5]), .ALUT(n13481[5]), .C0(n13490), 
          .Z(n13501[5]));
    LUT4 mux_4246_i2_3_lut (.A(dat_reg[9]), .B(dat_reg[1]), .C(n3980[4]), 
         .Z(n13481[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i2_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i2_3_lut (.A(dat_reg[25]), .B(dat_reg[17]), .C(n3980[2]), 
         .Z(n13471[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i2_3_lut.init = 16'hcaca;
    LUT4 mux_4246_i3_3_lut (.A(dat_reg[10]), .B(dat_reg[2]), .C(n3980[4]), 
         .Z(n13481[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i3_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i3_3_lut (.A(dat_reg[26]), .B(dat_reg[18]), .C(n3980[2]), 
         .Z(n13471[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i3_3_lut.init = 16'hcaca;
    LUT4 mux_4246_i4_3_lut (.A(dat_reg[11]), .B(dat_reg[3]), .C(n3980[4]), 
         .Z(n13481[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i4_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i4_3_lut (.A(dat_reg[27]), .B(dat_reg[19]), .C(n3980[2]), 
         .Z(n13471[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i4_3_lut.init = 16'hcaca;
    LUT4 mux_4246_i5_3_lut (.A(dat_reg[12]), .B(dat_reg[4]), .C(n3980[4]), 
         .Z(n13481[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i5_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i5_3_lut (.A(dat_reg[28]), .B(dat_reg[20]), .C(n3980[2]), 
         .Z(n13471[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i5_3_lut.init = 16'hcaca;
    LUT4 mux_4246_i6_3_lut (.A(dat_reg[13]), .B(dat_reg[5]), .C(n3980[4]), 
         .Z(n13481[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i6_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i6_3_lut (.A(dat_reg[29]), .B(dat_reg[21]), .C(n3980[2]), 
         .Z(n13471[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i6_3_lut.init = 16'hcaca;
    LUT4 mux_4246_i7_3_lut (.A(dat_reg[14]), .B(dat_reg[6]), .C(n3980[4]), 
         .Z(n13481[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i7_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i7_3_lut (.A(dat_reg[30]), .B(dat_reg[22]), .C(n3980[2]), 
         .Z(n13471[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i7_3_lut.init = 16'hcaca;
    PFUMX mux_4250_i5 (.BLUT(n13471[4]), .ALUT(n13481[4]), .C0(n13490), 
          .Z(n13501[4]));
    LUT4 i4248_2_lut (.A(n3980[3]), .B(n3980[4]), .Z(n13490)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i4248_2_lut.init = 16'heeee;
    LUT4 mux_4246_i8_3_lut (.A(dat_reg[15]), .B(dat_reg[7]), .C(n3980[4]), 
         .Z(n13481[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4246_i8_3_lut.init = 16'hcaca;
    LUT4 mux_4244_i8_3_lut (.A(dat_reg[31]), .B(dat_reg[23]), .C(n3980[2]), 
         .Z(n13471[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4244_i8_3_lut.init = 16'hcaca;
    PFUMX mux_4250_i4 (.BLUT(n13471[3]), .ALUT(n13481[3]), .C0(n13490), 
          .Z(n13501[3]));
    PFUMX mux_4250_i3 (.BLUT(n13471[2]), .ALUT(n13481[2]), .C0(n13490), 
          .Z(n13501[2]));
    PFUMX mux_4250_i2 (.BLUT(n13471[1]), .ALUT(n13481[1]), .C0(n13490), 
          .Z(n13501[1]));
    PFUMX mux_4250_i1 (.BLUT(n13471[0]), .ALUT(n13481[0]), .C0(n13490), 
          .Z(n13501[0]));
    
endmodule
//
// Verilog Description of module loadWeight
//

module loadWeight (sram_address_A, clock, n4445, sram_input_A, ramDataIn, 
            sram_ready_A, SDA_c, n73801, n1682, n1673, n73802, n39, 
            n23939, GND_net);
    output [11:0]sram_address_A;
    input clock;
    input n4445;
    output [31:0]sram_input_A;
    input [31:0]ramDataIn;
    output sram_ready_A;
    input SDA_c;
    input n73801;
    output n1682;
    output n1673;
    input n73802;
    input n39;
    input n23939;
    input GND_net;
    
    wire [31:0]addr;   // c:/users/yisong/documents/new/mlp/loadweight.vhd(40[8:12])
    wire n73801 /* synthesis nomerge= */ ;
    wire data_done;   // c:/users/yisong/documents/new/mlp/main.vhd(270[8:17])
    wire n73802 /* synthesis nomerge= */ ;
    
    wire n4810, n23636, n23863;
    wire [3:0]n1670;
    
    wire n30, n44, n38, n48, n34, n46, n52, n33, n42, n50, 
        n54, n41, n63345, n66251, n23683, n24027;
    wire [31:0]n134;
    
    wire n70722, n66534, n35176, n41_adj_569, n62727, n62726, n62725, 
        n62724, n62723, n62722, n62721, n62720, n62719, n62718, 
        n62717, n62716, n62715, n62714, n62713, n62712;
    
    FD1P3AX sram_addr_i0_i0 (.D(addr[0]), .SP(n4445), .CK(clock), .Q(sram_address_A[0]));
    defparam sram_addr_i0_i0.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i0 (.D(ramDataIn[0]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[0]));
    defparam sram_input_i0_i0.GSR = "DISABLED";
    FD1P3DX sram_ready_42 (.D(n23863), .SP(n23636), .CK(clock), .CD(SDA_c), 
            .Q(sram_ready_A));
    defparam sram_ready_42.GSR = "DISABLED";
    FD1S3BX state_FSM_i0 (.D(n73801), .CK(clock), .PD(SDA_c), .Q(n1670[0]));
    defparam state_FSM_i0.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i31 (.D(ramDataIn[31]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[31]));
    defparam sram_input_i0_i31.GSR = "DISABLED";
    LUT4 i2_2_lut (.A(addr[24]), .B(addr[1]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3AX sram_input_i0_i30 (.D(ramDataIn[30]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[30]));
    defparam sram_input_i0_i30.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i29 (.D(ramDataIn[29]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[29]));
    defparam sram_input_i0_i29.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i28 (.D(ramDataIn[28]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[28]));
    defparam sram_input_i0_i28.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i27 (.D(ramDataIn[27]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[27]));
    defparam sram_input_i0_i27.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i26 (.D(ramDataIn[26]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[26]));
    defparam sram_input_i0_i26.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i25 (.D(ramDataIn[25]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[25]));
    defparam sram_input_i0_i25.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i24 (.D(ramDataIn[24]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[24]));
    defparam sram_input_i0_i24.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i23 (.D(ramDataIn[23]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[23]));
    defparam sram_input_i0_i23.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i22 (.D(ramDataIn[22]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[22]));
    defparam sram_input_i0_i22.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i21 (.D(ramDataIn[21]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[21]));
    defparam sram_input_i0_i21.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i20 (.D(ramDataIn[20]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[20]));
    defparam sram_input_i0_i20.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i19 (.D(ramDataIn[19]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[19]));
    defparam sram_input_i0_i19.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i18 (.D(ramDataIn[18]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[18]));
    defparam sram_input_i0_i18.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i17 (.D(ramDataIn[17]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[17]));
    defparam sram_input_i0_i17.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i16 (.D(ramDataIn[16]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[16]));
    defparam sram_input_i0_i16.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i15 (.D(ramDataIn[15]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[15]));
    defparam sram_input_i0_i15.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i14 (.D(ramDataIn[14]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[14]));
    defparam sram_input_i0_i14.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i13 (.D(ramDataIn[13]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[13]));
    defparam sram_input_i0_i13.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i12 (.D(ramDataIn[12]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[12]));
    defparam sram_input_i0_i12.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i11 (.D(ramDataIn[11]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[11]));
    defparam sram_input_i0_i11.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i10 (.D(ramDataIn[10]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[10]));
    defparam sram_input_i0_i10.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i9 (.D(ramDataIn[9]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[9]));
    defparam sram_input_i0_i9.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i8 (.D(ramDataIn[8]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[8]));
    defparam sram_input_i0_i8.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i7 (.D(ramDataIn[7]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[7]));
    defparam sram_input_i0_i7.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i6 (.D(ramDataIn[6]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[6]));
    defparam sram_input_i0_i6.GSR = "DISABLED";
    LUT4 i16_4_lut (.A(addr[0]), .B(addr[7]), .C(addr[10]), .D(addr[15]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16_4_lut.init = 16'hfffe;
    FD1P3AX sram_input_i0_i5 (.D(ramDataIn[5]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[5]));
    defparam sram_input_i0_i5.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i4 (.D(ramDataIn[4]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[4]));
    defparam sram_input_i0_i4.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i3 (.D(ramDataIn[3]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[3]));
    defparam sram_input_i0_i3.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i2 (.D(ramDataIn[2]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[2]));
    defparam sram_input_i0_i2.GSR = "DISABLED";
    FD1P3AX sram_input_i0_i1 (.D(ramDataIn[1]), .SP(n4810), .CK(clock), 
            .Q(sram_input_A[1]));
    defparam sram_input_i0_i1.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i11 (.D(addr[11]), .SP(n4445), .CK(clock), .Q(sram_address_A[11]));
    defparam sram_addr_i0_i11.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i10 (.D(addr[10]), .SP(n4445), .CK(clock), .Q(sram_address_A[10]));
    defparam sram_addr_i0_i10.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i9 (.D(addr[9]), .SP(n4445), .CK(clock), .Q(sram_address_A[9]));
    defparam sram_addr_i0_i9.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i8 (.D(addr[8]), .SP(n4445), .CK(clock), .Q(sram_address_A[8]));
    defparam sram_addr_i0_i8.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i7 (.D(addr[7]), .SP(n4445), .CK(clock), .Q(sram_address_A[7]));
    defparam sram_addr_i0_i7.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i6 (.D(addr[6]), .SP(n4445), .CK(clock), .Q(sram_address_A[6]));
    defparam sram_addr_i0_i6.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i5 (.D(addr[5]), .SP(n4445), .CK(clock), .Q(sram_address_A[5]));
    defparam sram_addr_i0_i5.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i4 (.D(addr[4]), .SP(n4445), .CK(clock), .Q(sram_address_A[4]));
    defparam sram_addr_i0_i4.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i3 (.D(addr[3]), .SP(n4445), .CK(clock), .Q(sram_address_A[3]));
    defparam sram_addr_i0_i3.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i2 (.D(addr[2]), .SP(n4445), .CK(clock), .Q(sram_address_A[2]));
    defparam sram_addr_i0_i2.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i1 (.D(addr[1]), .SP(n4445), .CK(clock), .Q(sram_address_A[1]));
    defparam sram_addr_i0_i1.GSR = "DISABLED";
    LUT4 i10_2_lut (.A(addr[26]), .B(addr[6]), .Z(n38)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(addr[30]), .B(addr[13]), .C(addr[29]), .D(addr[28]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(addr[16]), .B(addr[9]), .Z(n34)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i18_4_lut (.A(addr[5]), .B(addr[27]), .C(addr[12]), .D(addr[14]), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(addr[11]), .B(n48), .C(n38), .D(addr[20]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(addr[18]), .B(addr[17]), .Z(n33)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i14_2_lut (.A(addr[19]), .B(addr[25]), .Z(n42)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(addr[8]), .B(n44), .C(n30), .D(addr[21]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(n33), .B(n52), .C(n46), .D(n34), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(addr[23]), .B(addr[22]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(n41), .B(n54), .C(n50), .D(n42), .Z(n63345)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut (.A(addr[3]), .B(addr[2]), .C(addr[31]), .D(addr[4]), 
         .Z(n66251)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i3_4_lut.init = 16'h0800;
    FD1P3IX addr_4651__i26 (.D(n134[26]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[26]));
    defparam addr_4651__i26.GSR = "DISABLED";
    FD1P3IX addr_4651__i29 (.D(n134[29]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[29]));
    defparam addr_4651__i29.GSR = "DISABLED";
    FD1P3IX addr_4651__i27 (.D(n134[27]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[27]));
    defparam addr_4651__i27.GSR = "DISABLED";
    FD1P3IX addr_4651__i30 (.D(n134[30]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[30]));
    defparam addr_4651__i30.GSR = "DISABLED";
    FD1P3IX addr_4651__i31 (.D(n134[31]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[31]));
    defparam addr_4651__i31.GSR = "DISABLED";
    FD1P3IX addr_4651__i28 (.D(n134[28]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[28]));
    defparam addr_4651__i28.GSR = "DISABLED";
    FD1P3IX addr_4651__i22 (.D(n134[22]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[22]));
    defparam addr_4651__i22.GSR = "DISABLED";
    FD1P3IX addr_4651__i16 (.D(n134[16]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[16]));
    defparam addr_4651__i16.GSR = "DISABLED";
    FD1P3IX addr_4651__i23 (.D(n134[23]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[23]));
    defparam addr_4651__i23.GSR = "DISABLED";
    FD1P3IX addr_4651__i17 (.D(n134[17]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[17]));
    defparam addr_4651__i17.GSR = "DISABLED";
    FD1P3IX addr_4651__i10 (.D(n134[10]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[10]));
    defparam addr_4651__i10.GSR = "DISABLED";
    FD1P3IX addr_4651__i12 (.D(n134[12]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[12]));
    defparam addr_4651__i12.GSR = "DISABLED";
    FD1P3IX addr_4651__i18 (.D(n134[18]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[18]));
    defparam addr_4651__i18.GSR = "DISABLED";
    FD1P3IX addr_4651__i24 (.D(n134[24]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[24]));
    defparam addr_4651__i24.GSR = "DISABLED";
    FD1P3IX addr_4651__i19 (.D(n134[19]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[19]));
    defparam addr_4651__i19.GSR = "DISABLED";
    FD1P3IX addr_4651__i13 (.D(n134[13]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[13]));
    defparam addr_4651__i13.GSR = "DISABLED";
    FD1P3IX addr_4651__i20 (.D(n134[20]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[20]));
    defparam addr_4651__i20.GSR = "DISABLED";
    FD1P3IX addr_4651__i14 (.D(n134[14]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[14]));
    defparam addr_4651__i14.GSR = "DISABLED";
    FD1P3IX addr_4651__i11 (.D(n134[11]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[11]));
    defparam addr_4651__i11.GSR = "DISABLED";
    FD1P3IX addr_4651__i15 (.D(n134[15]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[15]));
    defparam addr_4651__i15.GSR = "DISABLED";
    FD1P3IX addr_4651__i21 (.D(n134[21]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[21]));
    defparam addr_4651__i21.GSR = "DISABLED";
    FD1P3IX addr_4651__i25 (.D(n134[25]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[25]));
    defparam addr_4651__i25.GSR = "DISABLED";
    FD1P3IX addr_4651__i6 (.D(n134[6]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[6]));
    defparam addr_4651__i6.GSR = "DISABLED";
    FD1P3IX addr_4651__i7 (.D(n134[7]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[7]));
    defparam addr_4651__i7.GSR = "DISABLED";
    FD1P3IX addr_4651__i1 (.D(n134[1]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[1]));
    defparam addr_4651__i1.GSR = "DISABLED";
    FD1P3IX addr_4651__i2 (.D(n134[2]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[2]));
    defparam addr_4651__i2.GSR = "DISABLED";
    FD1P3IX addr_4651__i8 (.D(n134[8]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[8]));
    defparam addr_4651__i8.GSR = "DISABLED";
    FD1P3IX addr_4651__i3 (.D(n134[3]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[3]));
    defparam addr_4651__i3.GSR = "DISABLED";
    FD1P3IX addr_4651__i4 (.D(n134[4]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[4]));
    defparam addr_4651__i4.GSR = "DISABLED";
    FD1P3IX addr_4651__i5 (.D(n134[5]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[5]));
    defparam addr_4651__i5.GSR = "DISABLED";
    FD1P3IX addr_4651__i9 (.D(n134[9]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[9]));
    defparam addr_4651__i9.GSR = "DISABLED";
    LUT4 i12174_1_lut (.A(n1670[3]), .Z(n23863)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12174_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(n1670[0]), .B(n1670[3]), .Z(n23636)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i55095_3_lut_4_lut (.A(n66251), .B(n63345), .C(n1670[2]), .D(n23683), 
         .Z(n24027)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (C+!(D)))) */ ;
    defparam i55095_3_lut_4_lut.init = 16'h2f00;
    LUT4 i199_2_lut_3_lut (.A(n66251), .B(n63345), .C(n1670[2]), .Z(n1682)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i199_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_752 (.A(n66251), .B(n63345), .Z(n70722)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_752.init = 16'hdddd;
    LUT4 i2_3_lut (.A(n1673), .B(SDA_c), .C(data_done), .Z(n4810)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_3_lut.init = 16'h2020;
    FD1S3DX state_FSM_i1 (.D(n66534), .CK(clock), .CD(SDA_c), .Q(n1673));
    defparam state_FSM_i1.GSR = "DISABLED";
    FD1S3DX state_FSM_i2 (.D(n35176), .CK(clock), .CD(SDA_c), .Q(n1670[2]));
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1P3DX state_FSM_i3 (.D(n73802), .SP(n1682), .CK(clock), .CD(SDA_c), 
            .Q(n1670[3]));
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1P3IX addr_4651__i0 (.D(n134[0]), .SP(n23683), .CD(n24027), .CK(clock), 
            .Q(addr[0]));
    defparam addr_4651__i0.GSR = "DISABLED";
    FD1P3DX done_72 (.D(n23939), .SP(n39), .CK(clock), .CD(SDA_c), .Q(data_done));
    defparam done_72.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_981 (.A(data_done), .B(n1673), .Z(n35176)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_981.init = 16'h8888;
    LUT4 i1_3_lut (.A(n1670[2]), .B(n63345), .C(n66251), .Z(n41_adj_569)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h7575;
    LUT4 i1_4_lut (.A(n1670[0]), .B(data_done), .C(n41_adj_569), .D(n1673), 
         .Z(n66534)) /* synthesis lut_function=(A+!(B (C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'hbfaf;
    LUT4 i55080_4_lut (.A(n1670[0]), .B(SDA_c), .C(n70722), .D(n1670[2]), 
         .Z(n23683)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i55080_4_lut.init = 16'h3022;
    CCU2D addr_4651_add_4_33 (.A0(addr[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62727), .S0(n134[31]));
    defparam addr_4651_add_4_33.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_33.INIT1 = 16'h0000;
    defparam addr_4651_add_4_33.INJECT1_0 = "NO";
    defparam addr_4651_add_4_33.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_31 (.A0(addr[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62726), .COUT(n62727), .S0(n134[29]), .S1(n134[30]));
    defparam addr_4651_add_4_31.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_31.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_31.INJECT1_0 = "NO";
    defparam addr_4651_add_4_31.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_29 (.A0(addr[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62725), .COUT(n62726), .S0(n134[27]), .S1(n134[28]));
    defparam addr_4651_add_4_29.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_29.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_29.INJECT1_0 = "NO";
    defparam addr_4651_add_4_29.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_27 (.A0(addr[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62724), .COUT(n62725), .S0(n134[25]), .S1(n134[26]));
    defparam addr_4651_add_4_27.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_27.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_27.INJECT1_0 = "NO";
    defparam addr_4651_add_4_27.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_25 (.A0(addr[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62723), .COUT(n62724), .S0(n134[23]), .S1(n134[24]));
    defparam addr_4651_add_4_25.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_25.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_25.INJECT1_0 = "NO";
    defparam addr_4651_add_4_25.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_23 (.A0(addr[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62722), .COUT(n62723), .S0(n134[21]), .S1(n134[22]));
    defparam addr_4651_add_4_23.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_23.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_23.INJECT1_0 = "NO";
    defparam addr_4651_add_4_23.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_21 (.A0(addr[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62721), .COUT(n62722), .S0(n134[19]), .S1(n134[20]));
    defparam addr_4651_add_4_21.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_21.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_21.INJECT1_0 = "NO";
    defparam addr_4651_add_4_21.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_19 (.A0(addr[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62720), .COUT(n62721), .S0(n134[17]), .S1(n134[18]));
    defparam addr_4651_add_4_19.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_19.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_19.INJECT1_0 = "NO";
    defparam addr_4651_add_4_19.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_17 (.A0(addr[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62719), .COUT(n62720), .S0(n134[15]), .S1(n134[16]));
    defparam addr_4651_add_4_17.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_17.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_17.INJECT1_0 = "NO";
    defparam addr_4651_add_4_17.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_15 (.A0(addr[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62718), .COUT(n62719), .S0(n134[13]), .S1(n134[14]));
    defparam addr_4651_add_4_15.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_15.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_15.INJECT1_0 = "NO";
    defparam addr_4651_add_4_15.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_13 (.A0(addr[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62717), .COUT(n62718), .S0(n134[11]), .S1(n134[12]));
    defparam addr_4651_add_4_13.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_13.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_13.INJECT1_0 = "NO";
    defparam addr_4651_add_4_13.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_11 (.A0(addr[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62716), .COUT(n62717), .S0(n134[9]), .S1(n134[10]));
    defparam addr_4651_add_4_11.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_11.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_11.INJECT1_0 = "NO";
    defparam addr_4651_add_4_11.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_9 (.A0(addr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62715), .COUT(n62716), .S0(n134[7]), .S1(n134[8]));
    defparam addr_4651_add_4_9.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_9.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_9.INJECT1_0 = "NO";
    defparam addr_4651_add_4_9.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_7 (.A0(addr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62714), .COUT(n62715), .S0(n134[5]), .S1(n134[6]));
    defparam addr_4651_add_4_7.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_7.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_7.INJECT1_0 = "NO";
    defparam addr_4651_add_4_7.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_5 (.A0(addr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62713), .COUT(n62714), .S0(n134[3]), .S1(n134[4]));
    defparam addr_4651_add_4_5.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_5.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_5.INJECT1_0 = "NO";
    defparam addr_4651_add_4_5.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_3 (.A0(addr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62712), .COUT(n62713), .S0(n134[1]), .S1(n134[2]));
    defparam addr_4651_add_4_3.INIT0 = 16'hfaaa;
    defparam addr_4651_add_4_3.INIT1 = 16'hfaaa;
    defparam addr_4651_add_4_3.INJECT1_0 = "NO";
    defparam addr_4651_add_4_3.INJECT1_1 = "NO";
    CCU2D addr_4651_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n62712), .S1(n134[0]));
    defparam addr_4651_add_4_1.INIT0 = 16'hF000;
    defparam addr_4651_add_4_1.INIT1 = 16'h0555;
    defparam addr_4651_add_4_1.INJECT1_0 = "NO";
    defparam addr_4651_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module receiver
//

module receiver (clock, SDA_c, read_data, ramDataIn, count, n63477, 
            new_data, n25, n70855, GND_net);
    input clock;
    input SDA_c;
    input [7:0]read_data;
    output [31:0]ramDataIn;
    output [31:0]count;
    output n63477;
    input new_data;
    output n25;
    input n70855;
    input GND_net;
    
    wire [31:0]dat_reg;   // c:/users/yisong/documents/new/mlp/receiver.vhd(23[8:15])
    wire [31:0]count_c;   // c:/users/yisong/documents/new/mlp/receiver.vhd(20[8:13])
    
    wire n4438, n63, n19588, n19572, n19556;
    wire [31:0]n134;
    wire [31:0]n168;
    
    wire n70735, n32, n46, n40, n50, n36, n48, n54, n35, n44, 
        n52, n56, n43, n62743, n62742, n62741, n62740, n62739, 
        n62738, n62737, n62736, n62735, n62734, n62733, n62732, 
        n62731, n62730, n62729, n62728;
    
    FD1P3DX dat_reg_i0_i0 (.D(read_data[0]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[0]));
    defparam dat_reg_i0_i0.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i0 (.D(dat_reg[0]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[0]));
    defparam DataOut_i0_i0.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(count[1]), .B(count[0]), .C(count_c[2]), .D(n63477), 
         .Z(n63)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i3_4_lut.init = 16'hffef;
    LUT4 i8286_2_lut (.A(n63), .B(new_data), .Z(n19588)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i8286_2_lut.init = 16'h4444;
    FD1P3DX DataOut_i0_i31 (.D(dat_reg[31]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[31]));
    defparam DataOut_i0_i31.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i30 (.D(dat_reg[30]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[30]));
    defparam DataOut_i0_i30.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i29 (.D(dat_reg[29]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[29]));
    defparam DataOut_i0_i29.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i28 (.D(dat_reg[28]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[28]));
    defparam DataOut_i0_i28.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i27 (.D(dat_reg[27]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[27]));
    defparam DataOut_i0_i27.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i26 (.D(dat_reg[26]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[26]));
    defparam DataOut_i0_i26.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i25 (.D(dat_reg[25]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[25]));
    defparam DataOut_i0_i25.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i24 (.D(dat_reg[24]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[24]));
    defparam DataOut_i0_i24.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i23 (.D(dat_reg[23]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[23]));
    defparam DataOut_i0_i23.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i22 (.D(dat_reg[22]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[22]));
    defparam DataOut_i0_i22.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i21 (.D(dat_reg[21]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[21]));
    defparam DataOut_i0_i21.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i20 (.D(dat_reg[20]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[20]));
    defparam DataOut_i0_i20.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i19 (.D(dat_reg[19]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[19]));
    defparam DataOut_i0_i19.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i18 (.D(dat_reg[18]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[18]));
    defparam DataOut_i0_i18.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i17 (.D(dat_reg[17]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[17]));
    defparam DataOut_i0_i17.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i16 (.D(dat_reg[16]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[16]));
    defparam DataOut_i0_i16.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i15 (.D(dat_reg[15]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[15]));
    defparam DataOut_i0_i15.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i14 (.D(dat_reg[14]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[14]));
    defparam DataOut_i0_i14.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i13 (.D(dat_reg[13]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[13]));
    defparam DataOut_i0_i13.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i12 (.D(dat_reg[12]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[12]));
    defparam DataOut_i0_i12.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i11 (.D(dat_reg[11]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[11]));
    defparam DataOut_i0_i11.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i10 (.D(dat_reg[10]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[10]));
    defparam DataOut_i0_i10.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i9 (.D(dat_reg[9]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[9]));
    defparam DataOut_i0_i9.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i8 (.D(dat_reg[8]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[8]));
    defparam DataOut_i0_i8.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i7 (.D(dat_reg[7]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[7]));
    defparam DataOut_i0_i7.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i6 (.D(dat_reg[6]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[6]));
    defparam DataOut_i0_i6.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i5 (.D(dat_reg[5]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[5]));
    defparam DataOut_i0_i5.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i4 (.D(dat_reg[4]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[4]));
    defparam DataOut_i0_i4.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i3 (.D(dat_reg[3]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[3]));
    defparam DataOut_i0_i3.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i2 (.D(dat_reg[2]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[2]));
    defparam DataOut_i0_i2.GSR = "DISABLED";
    FD1P3DX DataOut_i0_i1 (.D(dat_reg[1]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(ramDataIn[1]));
    defparam DataOut_i0_i1.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i31 (.D(read_data[7]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[31]));
    defparam dat_reg_i0_i31.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i30 (.D(read_data[6]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[30]));
    defparam dat_reg_i0_i30.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i29 (.D(read_data[5]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[29]));
    defparam dat_reg_i0_i29.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i28 (.D(read_data[4]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[28]));
    defparam dat_reg_i0_i28.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i27 (.D(read_data[3]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[27]));
    defparam dat_reg_i0_i27.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i26 (.D(read_data[2]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[26]));
    defparam dat_reg_i0_i26.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i25 (.D(read_data[1]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[25]));
    defparam dat_reg_i0_i25.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i24 (.D(read_data[0]), .SP(n19588), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[24]));
    defparam dat_reg_i0_i24.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i23 (.D(read_data[7]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[23]));
    defparam dat_reg_i0_i23.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i22 (.D(read_data[6]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[22]));
    defparam dat_reg_i0_i22.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i21 (.D(read_data[5]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[21]));
    defparam dat_reg_i0_i21.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i20 (.D(read_data[4]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[20]));
    defparam dat_reg_i0_i20.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i19 (.D(read_data[3]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[19]));
    defparam dat_reg_i0_i19.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i18 (.D(read_data[2]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[18]));
    defparam dat_reg_i0_i18.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i17 (.D(read_data[1]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[17]));
    defparam dat_reg_i0_i17.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i16 (.D(read_data[0]), .SP(n19572), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[16]));
    defparam dat_reg_i0_i16.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i15 (.D(read_data[7]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[15]));
    defparam dat_reg_i0_i15.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i14 (.D(read_data[6]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[14]));
    defparam dat_reg_i0_i14.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i13 (.D(read_data[5]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[13]));
    defparam dat_reg_i0_i13.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i12 (.D(read_data[4]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[12]));
    defparam dat_reg_i0_i12.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i11 (.D(read_data[3]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[11]));
    defparam dat_reg_i0_i11.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i10 (.D(read_data[2]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[10]));
    defparam dat_reg_i0_i10.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i9 (.D(read_data[1]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[9]));
    defparam dat_reg_i0_i9.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i8 (.D(read_data[0]), .SP(n19556), .CK(clock), 
            .CD(SDA_c), .Q(dat_reg[8]));
    defparam dat_reg_i0_i8.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i7 (.D(read_data[7]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[7]));
    defparam dat_reg_i0_i7.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i6 (.D(read_data[6]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[6]));
    defparam dat_reg_i0_i6.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i5 (.D(read_data[5]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[5]));
    defparam dat_reg_i0_i5.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i4 (.D(read_data[4]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[4]));
    defparam dat_reg_i0_i4.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i3 (.D(read_data[3]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[3]));
    defparam dat_reg_i0_i3.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i2 (.D(read_data[2]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[2]));
    defparam dat_reg_i0_i2.GSR = "DISABLED";
    FD1P3DX dat_reg_i0_i1 (.D(read_data[1]), .SP(n4438), .CK(clock), .CD(SDA_c), 
            .Q(dat_reg[1]));
    defparam dat_reg_i0_i1.GSR = "DISABLED";
    LUT4 i34040_3_lut (.A(count[0]), .B(count_c[2]), .C(count[1]), .Z(n25)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i34040_3_lut.init = 16'hc9c9;
    LUT4 i29255_2_lut (.A(n134[31]), .B(n63), .Z(n168[31])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29255_2_lut.init = 16'h8888;
    LUT4 i29254_2_lut (.A(n134[30]), .B(n63), .Z(n168[30])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29254_2_lut.init = 16'h8888;
    LUT4 i29253_2_lut (.A(n134[29]), .B(n63), .Z(n168[29])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29253_2_lut.init = 16'h8888;
    LUT4 i29252_2_lut (.A(n134[28]), .B(n63), .Z(n168[28])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29252_2_lut.init = 16'h8888;
    LUT4 i29251_2_lut (.A(n134[27]), .B(n63), .Z(n168[27])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29251_2_lut.init = 16'h8888;
    LUT4 i29250_2_lut (.A(n134[26]), .B(n63), .Z(n168[26])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29250_2_lut.init = 16'h8888;
    LUT4 i29249_2_lut (.A(n134[25]), .B(n63), .Z(n168[25])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29249_2_lut.init = 16'h8888;
    LUT4 i29248_2_lut (.A(n134[24]), .B(n63), .Z(n168[24])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29248_2_lut.init = 16'h8888;
    LUT4 i29247_2_lut (.A(n134[23]), .B(n63), .Z(n168[23])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29247_2_lut.init = 16'h8888;
    LUT4 i29246_2_lut (.A(n134[22]), .B(n63), .Z(n168[22])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29246_2_lut.init = 16'h8888;
    LUT4 i29245_2_lut (.A(n134[21]), .B(n63), .Z(n168[21])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29245_2_lut.init = 16'h8888;
    LUT4 i29244_2_lut (.A(n134[20]), .B(n63), .Z(n168[20])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29244_2_lut.init = 16'h8888;
    LUT4 i29243_2_lut (.A(n134[19]), .B(n63), .Z(n168[19])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29243_2_lut.init = 16'h8888;
    LUT4 i29242_2_lut (.A(n134[18]), .B(n63), .Z(n168[18])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29242_2_lut.init = 16'h8888;
    LUT4 i29241_2_lut (.A(n134[17]), .B(n63), .Z(n168[17])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29241_2_lut.init = 16'h8888;
    LUT4 i29240_2_lut (.A(n134[16]), .B(n63), .Z(n168[16])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29240_2_lut.init = 16'h8888;
    LUT4 i29239_2_lut (.A(n134[15]), .B(n63), .Z(n168[15])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29239_2_lut.init = 16'h8888;
    LUT4 i29238_2_lut (.A(n134[14]), .B(n63), .Z(n168[14])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29238_2_lut.init = 16'h8888;
    LUT4 i29237_2_lut (.A(n134[13]), .B(n63), .Z(n168[13])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29237_2_lut.init = 16'h8888;
    LUT4 i29236_2_lut (.A(n134[12]), .B(n63), .Z(n168[12])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29236_2_lut.init = 16'h8888;
    LUT4 i29235_2_lut (.A(n134[11]), .B(n63), .Z(n168[11])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29235_2_lut.init = 16'h8888;
    LUT4 i29234_2_lut (.A(n134[10]), .B(n63), .Z(n168[10])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29234_2_lut.init = 16'h8888;
    LUT4 i29233_2_lut (.A(n134[9]), .B(n63), .Z(n168[9])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29233_2_lut.init = 16'h8888;
    LUT4 i29232_2_lut (.A(n134[8]), .B(n63), .Z(n168[8])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29232_2_lut.init = 16'h8888;
    LUT4 i29231_2_lut (.A(n134[7]), .B(n63), .Z(n168[7])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29231_2_lut.init = 16'h8888;
    LUT4 i29230_2_lut (.A(n134[6]), .B(n63), .Z(n168[6])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29230_2_lut.init = 16'h8888;
    LUT4 i29229_2_lut (.A(n134[5]), .B(n63), .Z(n168[5])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29229_2_lut.init = 16'h8888;
    LUT4 i29228_2_lut (.A(n134[4]), .B(n63), .Z(n168[4])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29228_2_lut.init = 16'h8888;
    LUT4 i29227_2_lut (.A(n134[3]), .B(n63), .Z(n168[3])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29227_2_lut.init = 16'h8888;
    LUT4 i29226_2_lut (.A(n134[2]), .B(n63), .Z(n168[2])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29226_2_lut.init = 16'h8888;
    LUT4 i29225_2_lut (.A(n134[1]), .B(n63), .Z(n168[1])) /* synthesis lut_function=(A (B)) */ ;
    defparam i29225_2_lut.init = 16'h8888;
    FD1S3DX count_4648__i0 (.D(n168[0]), .CK(new_data), .CD(SDA_c), .Q(count[0]));
    defparam count_4648__i0.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut (.A(count_c[2]), .B(n63477), .C(count[1]), .D(n70855), 
         .Z(n4438)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count_c[2]), .B(n63477), .C(n70855), 
         .D(count[1]), .Z(n19572)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_765 (.A(count_c[2]), .B(n63477), .Z(n70735)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_765.init = 16'heeee;
    LUT4 i2_3_lut_4_lut_adj_980 (.A(count[1]), .B(n70735), .C(new_data), 
         .D(count[0]), .Z(n19556)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_980.init = 16'h0020;
    LUT4 i3_2_lut (.A(count_c[29]), .B(count_c[19]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(count_c[10]), .B(count_c[7]), .C(count_c[11]), 
         .D(count_c[30]), .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i11_2_lut (.A(count_c[27]), .B(count_c[18]), .Z(n40)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11_2_lut.init = 16'heeee;
    LUT4 i21_4_lut (.A(count_c[16]), .B(count_c[23]), .C(count_c[31]), 
         .D(count_c[26]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i7_2_lut (.A(count_c[13]), .B(count_c[15]), .Z(n36)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(count_c[8]), .B(count_c[9]), .C(count_c[20]), .D(count_c[14]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i25_4_lut (.A(count_c[4]), .B(n50), .C(n40), .D(count_c[17]), 
         .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(count_c[6]), .B(count_c[12]), .Z(n35)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i15_3_lut (.A(count_c[28]), .B(count_c[22]), .C(count_c[25]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i23_4_lut (.A(count_c[3]), .B(n46), .C(n32), .D(count_c[5]), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i27_4_lut (.A(n35), .B(n54), .C(n48), .D(n36), .Z(n56)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut (.A(count_c[21]), .B(count_c[24]), .Z(n43)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i28_4_lut (.A(n43), .B(n56), .C(n52), .D(n44), .Z(n63477)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    FD1S3DX count_4648__i1 (.D(n168[1]), .CK(new_data), .CD(SDA_c), .Q(count[1]));
    defparam count_4648__i1.GSR = "DISABLED";
    FD1S3DX count_4648__i2 (.D(n168[2]), .CK(new_data), .CD(SDA_c), .Q(count_c[2]));
    defparam count_4648__i2.GSR = "DISABLED";
    FD1S3DX count_4648__i3 (.D(n168[3]), .CK(new_data), .CD(SDA_c), .Q(count_c[3]));
    defparam count_4648__i3.GSR = "DISABLED";
    FD1S3DX count_4648__i4 (.D(n168[4]), .CK(new_data), .CD(SDA_c), .Q(count_c[4]));
    defparam count_4648__i4.GSR = "DISABLED";
    FD1S3DX count_4648__i5 (.D(n168[5]), .CK(new_data), .CD(SDA_c), .Q(count_c[5]));
    defparam count_4648__i5.GSR = "DISABLED";
    FD1S3DX count_4648__i6 (.D(n168[6]), .CK(new_data), .CD(SDA_c), .Q(count_c[6]));
    defparam count_4648__i6.GSR = "DISABLED";
    FD1S3DX count_4648__i7 (.D(n168[7]), .CK(new_data), .CD(SDA_c), .Q(count_c[7]));
    defparam count_4648__i7.GSR = "DISABLED";
    FD1S3DX count_4648__i8 (.D(n168[8]), .CK(new_data), .CD(SDA_c), .Q(count_c[8]));
    defparam count_4648__i8.GSR = "DISABLED";
    FD1S3DX count_4648__i9 (.D(n168[9]), .CK(new_data), .CD(SDA_c), .Q(count_c[9]));
    defparam count_4648__i9.GSR = "DISABLED";
    FD1S3DX count_4648__i10 (.D(n168[10]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[10]));
    defparam count_4648__i10.GSR = "DISABLED";
    FD1S3DX count_4648__i11 (.D(n168[11]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[11]));
    defparam count_4648__i11.GSR = "DISABLED";
    FD1S3DX count_4648__i12 (.D(n168[12]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[12]));
    defparam count_4648__i12.GSR = "DISABLED";
    FD1S3DX count_4648__i13 (.D(n168[13]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[13]));
    defparam count_4648__i13.GSR = "DISABLED";
    FD1S3DX count_4648__i14 (.D(n168[14]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[14]));
    defparam count_4648__i14.GSR = "DISABLED";
    FD1S3DX count_4648__i15 (.D(n168[15]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[15]));
    defparam count_4648__i15.GSR = "DISABLED";
    FD1S3DX count_4648__i16 (.D(n168[16]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[16]));
    defparam count_4648__i16.GSR = "DISABLED";
    FD1S3DX count_4648__i17 (.D(n168[17]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[17]));
    defparam count_4648__i17.GSR = "DISABLED";
    FD1S3DX count_4648__i18 (.D(n168[18]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[18]));
    defparam count_4648__i18.GSR = "DISABLED";
    FD1S3DX count_4648__i19 (.D(n168[19]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[19]));
    defparam count_4648__i19.GSR = "DISABLED";
    FD1S3DX count_4648__i20 (.D(n168[20]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[20]));
    defparam count_4648__i20.GSR = "DISABLED";
    FD1S3DX count_4648__i21 (.D(n168[21]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[21]));
    defparam count_4648__i21.GSR = "DISABLED";
    FD1S3DX count_4648__i22 (.D(n168[22]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[22]));
    defparam count_4648__i22.GSR = "DISABLED";
    FD1S3DX count_4648__i23 (.D(n168[23]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[23]));
    defparam count_4648__i23.GSR = "DISABLED";
    FD1S3DX count_4648__i24 (.D(n168[24]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[24]));
    defparam count_4648__i24.GSR = "DISABLED";
    FD1S3DX count_4648__i25 (.D(n168[25]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[25]));
    defparam count_4648__i25.GSR = "DISABLED";
    FD1S3DX count_4648__i26 (.D(n168[26]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[26]));
    defparam count_4648__i26.GSR = "DISABLED";
    FD1S3DX count_4648__i27 (.D(n168[27]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[27]));
    defparam count_4648__i27.GSR = "DISABLED";
    FD1S3DX count_4648__i28 (.D(n168[28]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[28]));
    defparam count_4648__i28.GSR = "DISABLED";
    FD1S3DX count_4648__i29 (.D(n168[29]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[29]));
    defparam count_4648__i29.GSR = "DISABLED";
    FD1S3DX count_4648__i30 (.D(n168[30]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[30]));
    defparam count_4648__i30.GSR = "DISABLED";
    FD1S3DX count_4648__i31 (.D(n168[31]), .CK(new_data), .CD(SDA_c), 
            .Q(count_c[31]));
    defparam count_4648__i31.GSR = "DISABLED";
    LUT4 i28343_2_lut (.A(n134[0]), .B(n63), .Z(n168[0])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i28343_2_lut.init = 16'hbbbb;
    CCU2D count_4648_add_4_33 (.A0(count_c[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62743), .S0(n134[31]));
    defparam count_4648_add_4_33.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_33.INIT1 = 16'h0000;
    defparam count_4648_add_4_33.INJECT1_0 = "NO";
    defparam count_4648_add_4_33.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_31 (.A0(count_c[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62742), .COUT(n62743), .S0(n134[29]), 
          .S1(n134[30]));
    defparam count_4648_add_4_31.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_31.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_31.INJECT1_0 = "NO";
    defparam count_4648_add_4_31.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_29 (.A0(count_c[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62741), .COUT(n62742), .S0(n134[27]), 
          .S1(n134[28]));
    defparam count_4648_add_4_29.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_29.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_29.INJECT1_0 = "NO";
    defparam count_4648_add_4_29.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_27 (.A0(count_c[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62740), .COUT(n62741), .S0(n134[25]), 
          .S1(n134[26]));
    defparam count_4648_add_4_27.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_27.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_27.INJECT1_0 = "NO";
    defparam count_4648_add_4_27.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_25 (.A0(count_c[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62739), .COUT(n62740), .S0(n134[23]), 
          .S1(n134[24]));
    defparam count_4648_add_4_25.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_25.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_25.INJECT1_0 = "NO";
    defparam count_4648_add_4_25.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_23 (.A0(count_c[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62738), .COUT(n62739), .S0(n134[21]), 
          .S1(n134[22]));
    defparam count_4648_add_4_23.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_23.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_23.INJECT1_0 = "NO";
    defparam count_4648_add_4_23.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_21 (.A0(count_c[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62737), .COUT(n62738), .S0(n134[19]), 
          .S1(n134[20]));
    defparam count_4648_add_4_21.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_21.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_21.INJECT1_0 = "NO";
    defparam count_4648_add_4_21.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_19 (.A0(count_c[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62736), .COUT(n62737), .S0(n134[17]), 
          .S1(n134[18]));
    defparam count_4648_add_4_19.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_19.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_19.INJECT1_0 = "NO";
    defparam count_4648_add_4_19.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_17 (.A0(count_c[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62735), .COUT(n62736), .S0(n134[15]), 
          .S1(n134[16]));
    defparam count_4648_add_4_17.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_17.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_17.INJECT1_0 = "NO";
    defparam count_4648_add_4_17.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_15 (.A0(count_c[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62734), .COUT(n62735), .S0(n134[13]), 
          .S1(n134[14]));
    defparam count_4648_add_4_15.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_15.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_15.INJECT1_0 = "NO";
    defparam count_4648_add_4_15.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_13 (.A0(count_c[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62733), .COUT(n62734), .S0(n134[11]), 
          .S1(n134[12]));
    defparam count_4648_add_4_13.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_13.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_13.INJECT1_0 = "NO";
    defparam count_4648_add_4_13.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_11 (.A0(count_c[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62732), .COUT(n62733), .S0(n134[9]), .S1(n134[10]));
    defparam count_4648_add_4_11.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_11.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_11.INJECT1_0 = "NO";
    defparam count_4648_add_4_11.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_9 (.A0(count_c[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62731), .COUT(n62732), .S0(n134[7]), .S1(n134[8]));
    defparam count_4648_add_4_9.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_9.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_9.INJECT1_0 = "NO";
    defparam count_4648_add_4_9.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_7 (.A0(count_c[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62730), .COUT(n62731), .S0(n134[5]), .S1(n134[6]));
    defparam count_4648_add_4_7.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_7.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_7.INJECT1_0 = "NO";
    defparam count_4648_add_4_7.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_5 (.A0(count_c[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62729), .COUT(n62730), .S0(n134[3]), .S1(n134[4]));
    defparam count_4648_add_4_5.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_5.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_5.INJECT1_0 = "NO";
    defparam count_4648_add_4_5.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_3 (.A0(count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_c[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62728), .COUT(n62729), .S0(n134[1]), .S1(n134[2]));
    defparam count_4648_add_4_3.INIT0 = 16'hfaaa;
    defparam count_4648_add_4_3.INIT1 = 16'hfaaa;
    defparam count_4648_add_4_3.INJECT1_0 = "NO";
    defparam count_4648_add_4_3.INJECT1_1 = "NO";
    CCU2D count_4648_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n62728), .S1(n134[0]));
    defparam count_4648_add_4_1.INIT0 = 16'hF000;
    defparam count_4648_add_4_1.INIT1 = 16'h0555;
    defparam count_4648_add_4_1.INJECT1_0 = "NO";
    defparam count_4648_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module spi2
//

module spi2 (clock, new_data, GND_net, VCC_net, CE1_c, spi_mosi_oe, 
            spi_mosi_o, spi_miso_oe, spi_miso_o, spi_clk_oe, spi_clk_o, 
            spi_mosi_i, spi_miso_i, spi_clk_i, read_data, write_data, 
            n63477, n25, n39, \count[0] , \count[1] , n23939, n70855);
    input clock;
    output new_data;
    input GND_net;
    input VCC_net;
    input CE1_c;
    output spi_mosi_oe;
    output spi_mosi_o;
    output spi_miso_oe;
    output spi_miso_o;
    output spi_clk_oe;
    output spi_clk_o;
    input spi_mosi_i;
    input spi_miso_i;
    input spi_clk_i;
    output [7:0]read_data;
    input [7:0]write_data;
    input n63477;
    input n25;
    output n39;
    input \count[0] ;
    input \count[1] ;
    output n23939;
    output n70855;
    
    wire wbstb;   // c:/users/yisong/documents/new/mlp/spi.vhd(29[8:13])
    wire wback;   // c:/users/yisong/documents/new/mlp/spi.vhd(34[8:13])
    wire wbwe;   // c:/users/yisong/documents/new/mlp/spi.vhd(30[8:12])
    wire [7:0]wbaddr;   // c:/users/yisong/documents/new/mlp/spi.vhd(31[8:14])
    wire [7:0]wbdat_i;   // c:/users/yisong/documents/new/mlp/spi.vhd(32[8:15])
    wire [7:0]wbdat_o;   // c:/users/yisong/documents/new/mlp/spi.vhd(33[8:15])
    
    wire n40, n23823;
    wire [3:0]n1008;
    
    wire n70779, n17431, n70810, n29495, n32, n70811, n23645, 
        n47451, n70804, n35, n63303, n66103, n4637, n44;
    
    FD1S3IX wbstb_53 (.D(n40), .CK(clock), .CD(wback), .Q(wbstb));
    defparam wbstb_53.GSR = "DISABLED";
    FD1P3AX new_data_59 (.D(n1008[2]), .SP(n23823), .CK(clock), .Q(new_data));
    defparam new_data_59.GSR = "DISABLED";
    EFB EFBInst_0 (.WBCLKI(clock), .WBRSTI(GND_net), .WBCYCI(wbstb), .WBSTBI(wbstb), 
        .WBWEI(wbwe), .WBADRI0(wbaddr[0]), .WBADRI1(wbaddr[1]), .WBADRI2(wbaddr[2]), 
        .WBADRI3(wbaddr[3]), .WBADRI4(VCC_net), .WBADRI5(GND_net), .WBADRI6(VCC_net), 
        .WBADRI7(GND_net), .WBDATI0(wbdat_i[0]), .WBDATI1(wbdat_i[1]), 
        .WBDATI2(wbdat_i[2]), .WBDATI3(wbdat_i[3]), .WBDATI4(wbdat_i[4]), 
        .WBDATI5(wbdat_i[5]), .WBDATI6(wbdat_i[6]), .WBDATI7(wbdat_i[7]), 
        .I2C1SCLI(GND_net), .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), 
        .SPISCKI(spi_clk_i), .SPIMISOI(spi_miso_i), .SPIMOSII(spi_mosi_i), 
        .SPISCSN(CE1_c), .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), 
        .UFMSN(VCC_net), .PLL0DATI0(GND_net), .PLL0DATI1(GND_net), .PLL0DATI2(GND_net), 
        .PLL0DATI3(GND_net), .PLL0DATI4(GND_net), .PLL0DATI5(GND_net), 
        .PLL0DATI6(GND_net), .PLL0DATI7(GND_net), .PLL0ACKI(GND_net), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wbdat_o[0]), .WBDATO1(wbdat_o[1]), .WBDATO2(wbdat_o[2]), 
        .WBDATO3(wbdat_o[3]), .WBDATO4(wbdat_o[4]), .WBDATO5(wbdat_o[5]), 
        .WBDATO6(wbdat_o[6]), .WBDATO7(wbdat_o[7]), .WBACKO(wback), .SPISCKO(spi_clk_o), 
        .SPISCKEN(spi_clk_oe), .SPIMISOO(spi_miso_o), .SPIMISOEN(spi_miso_oe), 
        .SPIMOSIO(spi_mosi_o), .SPIMOSIEN(spi_mosi_oe)) /* synthesis syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/spi.vhd(48[8:27])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "ENABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "50.0";
    defparam EFBInst_0.DEV_DENSITY = "7000L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "SLAVE";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    FD1P3AX read_data_i0_i0 (.D(wbdat_o[0]), .SP(n70779), .CK(clock), 
            .Q(read_data[0]));
    defparam read_data_i0_i0.GSR = "DISABLED";
    FD1S3AX state_FSM_i1 (.D(n17431), .CK(clock), .Q(n1008[1]));
    defparam state_FSM_i1.GSR = "DISABLED";
    FD1P3AX wbaddr__i1 (.D(n29495), .SP(n70810), .CK(clock), .Q(wbaddr[0]));
    defparam wbaddr__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n1008[1]), .B(wbdat_o[4]), .C(n1008[3]), .D(wbdat_o[3]), 
         .Z(n32)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf0f2;
    LUT4 i1_2_lut_rep_841 (.A(n1008[1]), .B(wbdat_o[4]), .Z(n70811)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_841.init = 16'h2222;
    LUT4 i1_2_lut_2_lut (.A(wback), .B(n1008[3]), .Z(n23645)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i20_1_lut_rep_840 (.A(wback), .Z(n70810)) /* synthesis lut_function=(!(A)) */ ;
    defparam i20_1_lut_rep_840.init = 16'h5555;
    FD1P3IX wbdat_i_i0_i3 (.D(write_data[3]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[3]));
    defparam wbdat_i_i0_i3.GSR = "DISABLED";
    LUT4 i36110_1_lut_2_lut (.A(wback), .B(n1008[1]), .Z(n47451)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i36110_1_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_834 (.A(wback), .B(n1008[1]), .Z(n70804)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_834.init = 16'hbbbb;
    LUT4 i1_4_lut_4_lut (.A(wback), .B(n1008[2]), .C(n32), .D(n1008[1]), 
         .Z(n17431)) /* synthesis lut_function=(A (B+(C))+!A (D)) */ ;
    defparam i1_4_lut_4_lut.init = 16'hfda8;
    LUT4 i1_3_lut_3_lut (.A(wback), .B(n1008[2]), .C(n1008[1]), .Z(n23823)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam i1_3_lut_3_lut.init = 16'hb8b8;
    LUT4 i1_2_lut_rep_809 (.A(wback), .B(n1008[2]), .Z(n70779)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_809.init = 16'h8888;
    LUT4 i55128_2_lut (.A(n1008[1]), .B(n1008[2]), .Z(n35)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i55128_2_lut.init = 16'h1111;
    LUT4 i55083_3_lut (.A(new_data), .B(n63477), .C(n25), .Z(n39)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i55083_3_lut.init = 16'h5757;
    FD1P3IX wbdat_i_i0_i7 (.D(write_data[7]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[7]));
    defparam wbdat_i_i0_i7.GSR = "DISABLED";
    FD1S3JX state_FSM_i3 (.D(n63303), .CK(clock), .PD(n23645), .Q(n1008[3]));
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3AX state_FSM_i2 (.D(n66103), .CK(clock), .Q(n1008[2]));
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1P3AX read_data_i0_i7 (.D(wbdat_o[7]), .SP(n70779), .CK(clock), 
            .Q(read_data[7]));
    defparam read_data_i0_i7.GSR = "DISABLED";
    FD1P3AX read_data_i0_i6 (.D(wbdat_o[6]), .SP(n70779), .CK(clock), 
            .Q(read_data[6]));
    defparam read_data_i0_i6.GSR = "DISABLED";
    FD1P3AX read_data_i0_i5 (.D(wbdat_o[5]), .SP(n70779), .CK(clock), 
            .Q(read_data[5]));
    defparam read_data_i0_i5.GSR = "DISABLED";
    FD1P3AX read_data_i0_i4 (.D(wbdat_o[4]), .SP(n70779), .CK(clock), 
            .Q(read_data[4]));
    defparam read_data_i0_i4.GSR = "DISABLED";
    FD1P3AX read_data_i0_i3 (.D(wbdat_o[3]), .SP(n70779), .CK(clock), 
            .Q(read_data[3]));
    defparam read_data_i0_i3.GSR = "DISABLED";
    FD1P3AX read_data_i0_i2 (.D(wbdat_o[2]), .SP(n70779), .CK(clock), 
            .Q(read_data[2]));
    defparam read_data_i0_i2.GSR = "DISABLED";
    FD1P3AX read_data_i0_i1 (.D(wbdat_o[1]), .SP(n70779), .CK(clock), 
            .Q(read_data[1]));
    defparam read_data_i0_i1.GSR = "DISABLED";
    LUT4 i979_1_lut (.A(n1008[3]), .Z(n4637)) /* synthesis lut_function=(!(A)) */ ;
    defparam i979_1_lut.init = 16'h5555;
    FD1P3JX wbaddr__i2 (.D(n4637), .SP(n70810), .PD(n44), .CK(clock), 
            .Q(wbaddr[1]));
    defparam wbaddr__i2.GSR = "DISABLED";
    FD1P3IX wbaddr__i3 (.D(n70804), .SP(n70810), .CD(n29495), .CK(clock), 
            .Q(wbaddr[2]));
    defparam wbaddr__i3.GSR = "DISABLED";
    FD1P3JX wbaddr__i4 (.D(n47451), .SP(n70810), .PD(n29495), .CK(clock), 
            .Q(wbaddr[3]));
    defparam wbaddr__i4.GSR = "DISABLED";
    FD1P3IX wbdat_i_i0_i4 (.D(write_data[4]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[4]));
    defparam wbdat_i_i0_i4.GSR = "DISABLED";
    FD1P3IX wbdat_i_i0_i5 (.D(write_data[5]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[5]));
    defparam wbdat_i_i0_i5.GSR = "DISABLED";
    FD1P3IX wbdat_i_i0_i6 (.D(write_data[6]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[6]));
    defparam wbdat_i_i0_i6.GSR = "DISABLED";
    FD1S3IX wbwe_55 (.D(n35), .CK(clock), .CD(wback), .Q(wbwe));
    defparam wbwe_55.GSR = "DISABLED";
    FD1P3IX wbdat_i_i0_i0 (.D(write_data[0]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[0]));
    defparam wbdat_i_i0_i0.GSR = "DISABLED";
    FD1P3IX wbdat_i_i0_i1 (.D(write_data[1]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[1]));
    defparam wbdat_i_i0_i1.GSR = "DISABLED";
    FD1P3IX wbdat_i_i0_i2 (.D(write_data[2]), .SP(n23645), .CD(GND_net), 
            .CK(clock), .Q(wbdat_i[2]));
    defparam wbdat_i_i0_i2.GSR = "DISABLED";
    LUT4 i11_4_lut (.A(n1008[2]), .B(wbdat_o[3]), .C(wback), .D(n70811), 
         .Z(n66103)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i11_4_lut.init = 16'hca0a;
    LUT4 i2_3_lut (.A(wback), .B(wbdat_o[4]), .C(n1008[1]), .Z(n63303)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n1008[2]), .B(n1008[3]), .C(wback), 
         .Z(n29495)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i1_2_lut_3_lut (.A(n1008[2]), .B(n1008[3]), .C(n1008[1]), .Z(n40)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i55125_2_lut_2_lut_3_lut (.A(n1008[2]), .B(n1008[3]), .C(wback), 
         .Z(n44)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i55125_2_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_3_lut_adj_979 (.A(\count[0] ), .B(new_data), .C(\count[1] ), 
         .Z(n23939)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_979.init = 16'h0808;
    LUT4 i1_2_lut_rep_885 (.A(\count[0] ), .B(new_data), .Z(n70855)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_885.init = 16'h8888;
    
endmodule
//
// Verilog Description of module pr
//

module pr (n3946, clock, n23661, SDA_c, n73801, weight_done, n1682, 
           n73802, \state[0] , n3961, n3944, n22106);
    output n3946;
    input clock;
    input n23661;
    input SDA_c;
    input n73801;
    output weight_done;
    input n1682;
    input n73802;
    output \state[0] ;
    input n3961;
    output n3944;
    input n22106;
    
    wire n73801 /* synthesis nomerge= */ ;
    wire n73802 /* synthesis nomerge= */ ;
    
    FD1P3BX state_FSM__i1 (.D(n73801), .SP(n23661), .CK(clock), .PD(SDA_c), 
            .Q(n3946));
    defparam state_FSM__i1.GSR = "DISABLED";
    FD1P3DX weight_done_40 (.D(n73802), .SP(n1682), .CK(clock), .CD(SDA_c), 
            .Q(weight_done));
    defparam weight_done_40.GSR = "DISABLED";
    FD1P3DX state_FSM__i2 (.D(n3961), .SP(n23661), .CK(clock), .CD(SDA_c), 
            .Q(\state[0] ));
    defparam state_FSM__i2.GSR = "DISABLED";
    FD1P3DX state_FSM__i3 (.D(n22106), .SP(n23661), .CK(clock), .CD(SDA_c), 
            .Q(n3944));
    defparam state_FSM__i3.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module float_alu
//

module float_alu (n1151, n1156, \float_alu_mode[1] , \float_alu_mode[2] , 
            float_alu_c, clock, n70744, n70778, SDA_c, n70716, n24013, 
            n63113, n63130, float_alu_b, n62900, n124, float_alu_ready, 
            n70866, n2050, n4617, n2084, n15113, n2072, n4599, 
            n1155, n70822, n2036, n2086, n23655, n23979, n73809, 
            n70788, n73818, n2082, n23653, n45598, n63068, n62958, 
            n66522, n66524, n63156, n63069, n63070, n62961, n63102, 
            n63103, n63104, n63106, n63105, n63107, n63114, n63109, 
            n63115, n63116, n63120, n63122, n63128, n63131, n63139, 
            n63147, n63150, n62964, n62966, n1673, n4445, n27939, 
            n23942, n63112, n63111, n70816, GND_net, n42934, n61, 
            \A_int[10] , \B_int[10] , n70727, \A_int[11] , \B_int[11] , 
            \A_int[12] , \B_int[12] , n70692, \frac[15] , n70693, 
            \diffExpAB[8] , n493, n466, n70691, \efectFracB[13] , 
            \efectFracB[15] , \efectFracB[14] , \B_int[12]_adj_2 , \B_int[13] , 
            \B_int[15] , \B_int[8] , \A_int[2] , \A_int[3] , \A_int[6] , 
            \A_int[7] , \A_int[4] , \A_int[5] , \B_int[0] , \A_int[0] , 
            \A_int[11]_adj_3 , \A_int[12]_adj_4 , \A_int[13] , \A_int[15] , 
            \A_int[17] , \A_int[16] , \A_int[18] , \A_int[19] , \A_int[14] , 
            n4, n41520, \A_int[1] , \A_int[10]_adj_5 , \A_int[9] , 
            \A_int[22] , \A_int[21] , \A_int[8] , \A_int[20] , n22310, 
            \B_int[11]_adj_6 , \B_int[14] , \B_int[10]_adj_7 , \B_int[9] , 
            \B_int[19] , \B_int[18] , \B_int[20] , \B_int[21] , \B_int[7] , 
            n22437, \prod[47] , n66955, n67025, n67007, \prod[45] , 
            \prod[46] , \prod[28] , \prod[33] , \prod[40] , \prod[22] , 
            \prod[24] , \prod[25] , \prod[23] , \prod[26] , \prod[41] , 
            \prod[34] , \prod[37] , \prod[27] , \prod[39] , \prod[29] , 
            \prod[35] , \prod[36] , \prod[31] , \prod[32] , \prod[43] , 
            \prod[30] , \prod[38] , \prod[42] , \prod[44] , n42939, 
            n25571, \frac_norm[20] , \frac_norm[16] , \frac_norm[14] , 
            \frac_norm[15] , \frac_norm[12] , \frac_norm[13] , \frac_norm[10] , 
            \frac_norm[11] , \frac_norm[8] , n15, \B_int[17] , \B_int[16] , 
            \B_int[22] , \frac_norm[7] , n984, \B_int[3] , \B_int[1] , 
            \B_int[2] , \frac_norm[4] , \frac_norm[5] , \frac_norm[3] , 
            \frac_norm[2] , exp_final, \FP_Z_int[22] , \B_int[6] , \B_int[5] , 
            \B_int[4] , n6, \prod[21] , VCC_net, \buf_x[89] , \buf_x[87] , 
            \buf_x[88] , \buf_x[85] , \buf_x[86] , \buf_x[83] , \buf_x[84] , 
            \buf_r[89] , \buf_r[87] , \buf_r[88] , \buf_r[85] , \buf_r[86] , 
            \buf_r[83] , \buf_r[84] , \A_int[11]_adj_8 , \B_int[11]_adj_9 , 
            \A_int[10]_adj_10 , \B_int[10]_adj_11 , \A_int[13]_adj_12 , 
            \B_int[13]_adj_13 , \A_int[12]_adj_14 , \B_int[12]_adj_15 , 
            \A_int[17]_adj_16 , \B_int[17]_adj_17 , \A_int[16]_adj_18 , 
            \B_int[16]_adj_19 , \A_int[18]_adj_20 , \B_int[18]_adj_21 , 
            \A_int[2]_adj_22 , \B_int[2]_adj_23 , \B_int[3]_adj_24 , \A_int[9]_adj_25 , 
            \A_int[7]_adj_26 , \A_int[4]_adj_27 , \A_int[3]_adj_28 , \B_int[9]_adj_29 , 
            \B_int[7]_adj_30 , \B_int[4]_adj_31 , \diffExpAB[8]_adj_32 , 
            \diffExp[4] , n70835, n70834, n70833, \efectFracB[21] , 
            \efectFracB[20] , \efectFracB[19] , \efectFracB[15]_adj_33 , 
            \efectFracB[16] , n19214, n28, n70771, n9, \efectFracB[14]_adj_34 , 
            \efectFracB[7] , \efectFracB[5] , \efectFracB[12] , n70820, 
            \efectFracB[13]_adj_35 , n27, n70740, n55);
    output n1151;
    output n1156;
    input \float_alu_mode[1] ;
    input \float_alu_mode[2] ;
    output [31:0]float_alu_c;
    input clock;
    input n70744;
    output n70778;
    input SDA_c;
    input n70716;
    input n24013;
    input n63113;
    input n63130;
    input [31:0]float_alu_b;
    input n62900;
    input n124;
    input float_alu_ready;
    output n70866;
    input n2050;
    output n4617;
    input n2084;
    output n15113;
    input n2072;
    output n4599;
    output n1155;
    output n70822;
    input n2036;
    input n2086;
    output n23655;
    input n23979;
    output n73809;
    output n70788;
    output n73818;
    input n2082;
    output n23653;
    input n45598;
    input n63068;
    input n62958;
    input n66522;
    input n66524;
    input n63156;
    input n63069;
    input n63070;
    input n62961;
    input n63102;
    input n63103;
    input n63104;
    input n63106;
    input n63105;
    input n63107;
    input n63114;
    input n63109;
    input n63115;
    input n63116;
    input n63120;
    input n63122;
    input n63128;
    input n63131;
    input n63139;
    input n63147;
    input n63150;
    input n62964;
    input n62966;
    input n1673;
    output n4445;
    input n27939;
    input n23942;
    input n63112;
    input n63111;
    output n70816;
    input GND_net;
    input n42934;
    output n61;
    output \A_int[10] ;
    output \B_int[10] ;
    output n70727;
    output \A_int[11] ;
    output \B_int[11] ;
    output \A_int[12] ;
    output \B_int[12] ;
    input n70692;
    input \frac[15] ;
    output n70693;
    output \diffExpAB[8] ;
    output n493;
    output n466;
    input n70691;
    input \efectFracB[13] ;
    input \efectFracB[15] ;
    input \efectFracB[14] ;
    output \B_int[12]_adj_2 ;
    output \B_int[13] ;
    output \B_int[15] ;
    output \B_int[8] ;
    output \A_int[2] ;
    output \A_int[3] ;
    output \A_int[6] ;
    output \A_int[7] ;
    output \A_int[4] ;
    output \A_int[5] ;
    output \B_int[0] ;
    output \A_int[0] ;
    output \A_int[11]_adj_3 ;
    output \A_int[12]_adj_4 ;
    output \A_int[13] ;
    output \A_int[15] ;
    output \A_int[17] ;
    output \A_int[16] ;
    output \A_int[18] ;
    output \A_int[19] ;
    output \A_int[14] ;
    output n4;
    output n41520;
    output \A_int[1] ;
    output \A_int[10]_adj_5 ;
    output \A_int[9] ;
    output \A_int[22] ;
    output \A_int[21] ;
    output \A_int[8] ;
    output \A_int[20] ;
    output n22310;
    output \B_int[11]_adj_6 ;
    output \B_int[14] ;
    output \B_int[10]_adj_7 ;
    output \B_int[9] ;
    output \B_int[19] ;
    output \B_int[18] ;
    output \B_int[20] ;
    output \B_int[21] ;
    output \B_int[7] ;
    output n22437;
    input \prod[47] ;
    input n66955;
    input n67025;
    input n67007;
    input \prod[45] ;
    input \prod[46] ;
    input \prod[28] ;
    input \prod[33] ;
    input \prod[40] ;
    input \prod[22] ;
    input \prod[24] ;
    input \prod[25] ;
    input \prod[23] ;
    input \prod[26] ;
    input \prod[41] ;
    input \prod[34] ;
    input \prod[37] ;
    input \prod[27] ;
    input \prod[39] ;
    input \prod[29] ;
    input \prod[35] ;
    input \prod[36] ;
    input \prod[31] ;
    input \prod[32] ;
    input \prod[43] ;
    input \prod[30] ;
    input \prod[38] ;
    input \prod[42] ;
    input \prod[44] ;
    output n42939;
    output n25571;
    input \frac_norm[20] ;
    input \frac_norm[16] ;
    input \frac_norm[14] ;
    input \frac_norm[15] ;
    input \frac_norm[12] ;
    input \frac_norm[13] ;
    input \frac_norm[10] ;
    input \frac_norm[11] ;
    input \frac_norm[8] ;
    input n15;
    output \B_int[17] ;
    output \B_int[16] ;
    output \B_int[22] ;
    input \frac_norm[7] ;
    input [7:0]n984;
    output \B_int[3] ;
    output \B_int[1] ;
    output \B_int[2] ;
    input \frac_norm[4] ;
    input \frac_norm[5] ;
    input \frac_norm[3] ;
    input \frac_norm[2] ;
    output [7:0]exp_final;
    input \FP_Z_int[22] ;
    output \B_int[6] ;
    output \B_int[5] ;
    output \B_int[4] ;
    output n6;
    input \prod[21] ;
    input VCC_net;
    output \buf_x[89] ;
    output \buf_x[87] ;
    output \buf_x[88] ;
    output \buf_x[85] ;
    output \buf_x[86] ;
    output \buf_x[83] ;
    output \buf_x[84] ;
    input \buf_r[89] ;
    input \buf_r[87] ;
    input \buf_r[88] ;
    input \buf_r[85] ;
    input \buf_r[86] ;
    input \buf_r[83] ;
    input \buf_r[84] ;
    output \A_int[11]_adj_8 ;
    output \B_int[11]_adj_9 ;
    output \A_int[10]_adj_10 ;
    output \B_int[10]_adj_11 ;
    output \A_int[13]_adj_12 ;
    output \B_int[13]_adj_13 ;
    output \A_int[12]_adj_14 ;
    output \B_int[12]_adj_15 ;
    output \A_int[17]_adj_16 ;
    output \B_int[17]_adj_17 ;
    output \A_int[16]_adj_18 ;
    output \B_int[16]_adj_19 ;
    output \A_int[18]_adj_20 ;
    output \B_int[18]_adj_21 ;
    output \A_int[2]_adj_22 ;
    output \B_int[2]_adj_23 ;
    output \B_int[3]_adj_24 ;
    output \A_int[9]_adj_25 ;
    output \A_int[7]_adj_26 ;
    output \A_int[4]_adj_27 ;
    output \A_int[3]_adj_28 ;
    output \B_int[9]_adj_29 ;
    output \B_int[7]_adj_30 ;
    output \B_int[4]_adj_31 ;
    output \diffExpAB[8]_adj_32 ;
    output \diffExp[4] ;
    output n70835;
    output n70834;
    output n70833;
    input \efectFracB[21] ;
    input \efectFracB[20] ;
    input \efectFracB[19] ;
    input \efectFracB[15]_adj_33 ;
    input \efectFracB[16] ;
    input n19214;
    input n28;
    input n70771;
    input n9;
    input \efectFracB[14]_adj_34 ;
    input \efectFracB[7] ;
    input \efectFracB[5] ;
    input \efectFracB[12] ;
    input n70820;
    input \efectFracB[13]_adj_35 ;
    input n27;
    input n70740;
    input n55;
    
    wire [23:0]fR1_e3;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(820[10:16])
    wire ufl1_e3;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(831[10:17])
    wire [2:0]float_alu_mode;   // c:/users/yisong/documents/new/mlp/main.vhd(298[8:22])
    wire [31:0]wait_counter;   // c:/users/yisong/documents/new/mlp/fp.vhd(141[8:20])
    wire [31:0]add_c;   // c:/users/yisong/documents/new/mlp/fp.vhd(151[29:34])
    wire [31:0]sub_c;   // c:/users/yisong/documents/new/mlp/fp.vhd(151[36:41])
    wire [31:0]mul_c;   // c:/users/yisong/documents/new/mlp/fp.vhd(151[43:48])
    wire [31:0]div_c;   // c:/users/yisong/documents/new/mlp/fp.vhd(151[50:55])
    wire [31:0]float_alu_a;   // c:/users/yisong/documents/new/mlp/main.vhd(297[8:19])
    wire [31:0]alu_b;   // c:/users/yisong/documents/new/mlp/fp.vhd(151[15:20])
    wire add_ce;   // c:/users/yisong/documents/new/mlp/fp.vhd(145[8:14])
    wire sub_ce;   // c:/users/yisong/documents/new/mlp/fp.vhd(145[16:22])
    wire add_enable;   // c:/users/yisong/documents/new/mlp/fp.vhd(146[8:18])
    wire [31:0]alu_a;   // c:/users/yisong/documents/new/mlp/fp.vhd(151[8:13])
    wire [8:0]eR_e3;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(823[10:15])
    wire [24:0]mXs_0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(542[10:15])
    wire [33:0]exp_a;   // c:/users/yisong/documents/new/mlp/fp.vhd(148[8:13])
    wire mul_ce;   // c:/users/yisong/documents/new/mlp/fp.vhd(145[24:30])
    wire div_ce;   // c:/users/yisong/documents/new/mlp/fp.vhd(145[32:38])
    wire [31:0]n13301;
    wire [31:0]n13369;
    
    wire n22189, n24, n70814;
    wire [7:0]n1148;
    wire [31:0]n13267;
    
    wire n26, n20, n28_c;
    wire [31:0]n13437;
    
    wire n70781, n142, n47, n70841, n16, n66208, n10, n113, 
        n66700, n14, n73817, n73820, n23974, n23819, n67175, n70850, 
        n110, n23670, n23885, n66613, n23632, n45611, n142_adj_528, 
        n70790, n141, n70767;
    wire [30:0]n130;
    
    wire n23850, n23854, n23856, n23858, n23860, n23862, n23871, 
        n23877, n23882, n23884, n23891, n23893, n23895, n23897, 
        n23899, n23901, n23903, n23905, n23911, n23913, n23867, 
        n23873, n23917, n23919, n23921, n66808, n65745;
    wire [30:0]n163;
    
    wire n23915, n23875, n23722, n23972, n66655, n22185, n22187, 
        n70793, n45720, n16_adj_531, n17, n139_adj_532, n12, n4_c, 
        n66575, n73816, n69007, n70856, n1442, n68796, n86, n73804, 
        n70815, n73803, n69006, n70849, n68795, n62758, n62757, 
        n62756, n62755, n62754, n73815, n62753, n73812, n41808, 
        n42941, n25583, n62752, n62751, n62750, n62749, n62748, 
        n62747, n62746, n62745, n62744, n73814, n73813, n73811, 
        n73810;
    
    LUT4 i54891_4_lut (.A(n13301[3]), .B(fR1_e3[3]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54891_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1156), .B(float_alu_mode[0]), .C(\float_alu_mode[1] ), 
         .D(\float_alu_mode[2] ), .Z(n22189)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i9_4_lut (.A(wait_counter[4]), .B(wait_counter[18]), .C(wait_counter[9]), 
         .D(wait_counter[25]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_844_3_lut (.A(n1156), .B(float_alu_mode[0]), .C(\float_alu_mode[2] ), 
         .Z(n70814)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_844_3_lut.init = 16'h2020;
    LUT4 mux_4232_i4_3_lut (.A(add_c[3]), .B(sub_c[3]), .C(n1148[2]), 
         .Z(n13267[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i4_3_lut.init = 16'hcaca;
    LUT4 i13_4_lut (.A(wait_counter[6]), .B(n26), .C(n20), .D(wait_counter[14]), 
         .Z(n28_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 mux_4234_i5_3_lut (.A(mul_c[4]), .B(div_c[4]), .C(n1148[4]), 
         .Z(n13301[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i5_3_lut.init = 16'hcaca;
    LUT4 i54889_4_lut (.A(n13301[4]), .B(fR1_e3[4]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54889_4_lut.init = 16'h0aca;
    FD1P3AX alu_c_i0_i0 (.D(n13437[0]), .SP(n70744), .CK(clock), .Q(float_alu_c[0]));
    defparam alu_c_i0_i0.GSR = "DISABLED";
    LUT4 mux_4232_i5_3_lut (.A(add_c[4]), .B(sub_c[4]), .C(n1148[2]), 
         .Z(n13267[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i5_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_811_3_lut (.A(n1156), .B(float_alu_mode[0]), .C(\float_alu_mode[1] ), 
         .Z(n70781)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_811_3_lut.init = 16'h2020;
    LUT4 i129_3_lut_4_lut_3_lut (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .Z(n142)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;
    defparam i129_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 mux_4234_i6_3_lut (.A(mul_c[5]), .B(div_c[5]), .C(n1148[4]), 
         .Z(n13301[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i6_3_lut.init = 16'hcaca;
    LUT4 i54887_4_lut (.A(n13301[5]), .B(fR1_e3[5]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54887_4_lut.init = 16'h0aca;
    LUT4 i36_3_lut_4_lut_3_lut (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .Z(n47)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;
    defparam i36_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_4232_i6_3_lut (.A(add_c[5]), .B(sub_c[5]), .C(n1148[2]), 
         .Z(n13267[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i6_3_lut.init = 16'hcaca;
    LUT4 i2_1_lut_rep_871 (.A(\float_alu_mode[2] ), .Z(n70841)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut_rep_871.init = 16'h5555;
    LUT4 mux_4234_i7_3_lut (.A(mul_c[6]), .B(div_c[6]), .C(n1148[4]), 
         .Z(n13301[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i7_3_lut.init = 16'hcaca;
    LUT4 i54885_4_lut (.A(n13301[6]), .B(fR1_e3[6]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54885_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i7_3_lut (.A(add_c[6]), .B(sub_c[6]), .C(n1148[2]), 
         .Z(n13267[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i7_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i8_3_lut (.A(mul_c[7]), .B(div_c[7]), .C(n1148[4]), 
         .Z(n13301[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i8_3_lut.init = 16'hcaca;
    LUT4 i14_4_lut (.A(wait_counter[13]), .B(n28_c), .C(n24), .D(n16), 
         .Z(n66208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i54883_4_lut (.A(n13301[7]), .B(fR1_e3[7]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54883_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i8_3_lut (.A(add_c[7]), .B(sub_c[7]), .C(n1148[2]), 
         .Z(n13267[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i8_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i9_3_lut (.A(mul_c[8]), .B(div_c[8]), .C(n1148[4]), 
         .Z(n13301[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i9_3_lut.init = 16'hcaca;
    LUT4 i54881_4_lut (.A(n13301[8]), .B(fR1_e3[8]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54881_4_lut.init = 16'h0aca;
    LUT4 i2_2_lut (.A(wait_counter[22]), .B(wait_counter[20]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    FD1P3BX state_FSM__i1 (.D(n113), .SP(n70778), .CK(clock), .PD(SDA_c), 
            .Q(n1156));
    defparam state_FSM__i1.GSR = "DISABLED";
    LUT4 mux_4232_i9_3_lut (.A(add_c[8]), .B(sub_c[8]), .C(n1148[2]), 
         .Z(n13267[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i9_3_lut.init = 16'hcaca;
    LUT4 i6_4_lut (.A(wait_counter[24]), .B(wait_counter[23]), .C(n66208), 
         .D(n66700), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 mux_4234_i10_3_lut (.A(mul_c[9]), .B(div_c[9]), .C(n1148[4]), 
         .Z(n13301[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i10_3_lut.init = 16'hcaca;
    LUT4 i54879_4_lut (.A(n13301[9]), .B(fR1_e3[9]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54879_4_lut.init = 16'h0aca;
    FD1P3JX float_alu_a_i0_i28 (.D(n63113), .SP(n70716), .PD(n24013), 
            .CK(clock), .Q(float_alu_a[28]));
    defparam float_alu_a_i0_i28.GSR = "DISABLED";
    LUT4 mux_4232_i10_3_lut (.A(add_c[9]), .B(sub_c[9]), .C(n1148[2]), 
         .Z(n13267[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i10_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i11_3_lut (.A(mul_c[10]), .B(div_c[10]), .C(n1148[4]), 
         .Z(n13301[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i11_3_lut.init = 16'hcaca;
    LUT4 i54877_4_lut (.A(n13301[10]), .B(fR1_e3[10]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54877_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i11_3_lut (.A(add_c[10]), .B(sub_c[10]), .C(n1148[2]), 
         .Z(n13267[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i11_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i12_3_lut (.A(mul_c[11]), .B(div_c[11]), .C(n1148[4]), 
         .Z(n13301[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i12_3_lut.init = 16'hcaca;
    LUT4 i54875_4_lut (.A(n13301[11]), .B(fR1_e3[11]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54875_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i12_3_lut (.A(add_c[11]), .B(sub_c[11]), .C(n1148[2]), 
         .Z(n13267[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i12_3_lut.init = 16'hcaca;
    FD1P3JX float_alu_a_i0_i29 (.D(n63130), .SP(n70716), .PD(n24013), 
            .CK(clock), .Q(float_alu_a[29]));
    defparam float_alu_a_i0_i29.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i1 (.D(float_alu_b[1]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[1]));
    defparam alu_b_i0_i1.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i2 (.D(float_alu_b[2]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[2]));
    defparam alu_b_i0_i2.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i3 (.D(float_alu_b[3]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[3]));
    defparam alu_b_i0_i3.GSR = "DISABLED";
    LUT4 mux_4234_i13_3_lut (.A(mul_c[12]), .B(div_c[12]), .C(n1148[4]), 
         .Z(n13301[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i13_3_lut.init = 16'hcaca;
    LUT4 i54873_4_lut (.A(n13301[12]), .B(fR1_e3[12]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54873_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i13_3_lut (.A(add_c[12]), .B(sub_c[12]), .C(n1148[2]), 
         .Z(n13267[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i13_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i14_3_lut (.A(mul_c[13]), .B(div_c[13]), .C(n1148[4]), 
         .Z(n13301[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i14_3_lut.init = 16'hcaca;
    LUT4 i54871_4_lut (.A(n13301[13]), .B(fR1_e3[13]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54871_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i14_3_lut (.A(add_c[13]), .B(sub_c[13]), .C(n1148[2]), 
         .Z(n13267[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i14_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i15_3_lut (.A(mul_c[14]), .B(div_c[14]), .C(n1148[4]), 
         .Z(n13301[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i15_3_lut.init = 16'hcaca;
    LUT4 i54869_4_lut (.A(n13301[14]), .B(fR1_e3[14]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54869_4_lut.init = 16'h0aca;
    FD1P3IX alu_b_i0_i4 (.D(float_alu_b[4]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[4]));
    defparam alu_b_i0_i4.GSR = "DISABLED";
    LUT4 mux_4232_i15_3_lut (.A(add_c[14]), .B(sub_c[14]), .C(n1148[2]), 
         .Z(n13267[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i15_3_lut.init = 16'hcaca;
    FD1P3AX float_alu_a_i0_i0 (.D(n62900), .SP(n70716), .CK(clock), .Q(float_alu_a[0]));
    defparam float_alu_a_i0_i0.GSR = "DISABLED";
    LUT4 mux_4234_i16_3_lut (.A(mul_c[15]), .B(div_c[15]), .C(n1148[4]), 
         .Z(n13301[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i16_3_lut.init = 16'hcaca;
    LUT4 i54867_4_lut (.A(n13301[15]), .B(fR1_e3[15]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54867_4_lut.init = 16'h0aca;
    FD1P3IX alu_b_i0_i5 (.D(float_alu_b[5]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[5]));
    defparam alu_b_i0_i5.GSR = "DISABLED";
    LUT4 mux_4232_i16_3_lut (.A(add_c[15]), .B(sub_c[15]), .C(n1148[2]), 
         .Z(n13267[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i16_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i17_3_lut (.A(mul_c[16]), .B(div_c[16]), .C(n1148[4]), 
         .Z(n13301[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i17_3_lut.init = 16'hcaca;
    LUT4 i54865_4_lut (.A(n13301[16]), .B(fR1_e3[16]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54865_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i17_3_lut (.A(add_c[16]), .B(sub_c[16]), .C(n1148[2]), 
         .Z(n13267[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i17_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i18_3_lut (.A(mul_c[17]), .B(div_c[17]), .C(n1148[4]), 
         .Z(n13301[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i18_3_lut.init = 16'hcaca;
    LUT4 i54863_4_lut (.A(n13301[17]), .B(fR1_e3[17]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54863_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i18_3_lut (.A(add_c[17]), .B(sub_c[17]), .C(n1148[2]), 
         .Z(n13267[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i18_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i19_3_lut (.A(mul_c[18]), .B(div_c[18]), .C(n1148[4]), 
         .Z(n13301[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i19_3_lut.init = 16'hcaca;
    LUT4 i54861_4_lut (.A(n13301[18]), .B(fR1_e3[18]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54861_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i19_3_lut (.A(add_c[18]), .B(sub_c[18]), .C(n1148[2]), 
         .Z(n13267[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i19_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i20_3_lut (.A(mul_c[19]), .B(div_c[19]), .C(n1148[4]), 
         .Z(n13301[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i20_3_lut.init = 16'hcaca;
    LUT4 i54859_4_lut (.A(n13301[19]), .B(fR1_e3[19]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54859_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i20_3_lut (.A(add_c[19]), .B(sub_c[19]), .C(n1148[2]), 
         .Z(n13267[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i20_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i21_3_lut (.A(mul_c[20]), .B(div_c[20]), .C(n1148[4]), 
         .Z(n13301[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i21_3_lut.init = 16'hcaca;
    LUT4 i54857_4_lut (.A(n13301[20]), .B(fR1_e3[20]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54857_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i21_3_lut (.A(add_c[20]), .B(sub_c[20]), .C(n1148[2]), 
         .Z(n13267[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i21_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i22_3_lut (.A(mul_c[21]), .B(div_c[21]), .C(n1148[4]), 
         .Z(n13301[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i22_3_lut.init = 16'hcaca;
    LUT4 i54855_4_lut (.A(n13301[21]), .B(fR1_e3[21]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54855_4_lut.init = 16'h0aca;
    FD1P3AX add_ce_79 (.D(n124), .SP(n23819), .CK(clock), .Q(add_ce));
    defparam add_ce_79.GSR = "DISABLED";
    LUT4 mux_4232_i22_3_lut (.A(add_c[21]), .B(sub_c[21]), .C(n1148[2]), 
         .Z(n13267[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i22_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i23_3_lut (.A(mul_c[22]), .B(div_c[22]), .C(n1148[4]), 
         .Z(n13301[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i23_3_lut.init = 16'hcaca;
    FD1P3IX alu_b_i0_i6 (.D(float_alu_b[6]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[6]));
    defparam alu_b_i0_i6.GSR = "DISABLED";
    LUT4 i54853_4_lut (.A(n13301[22]), .B(fR1_e3[22]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54853_4_lut.init = 16'h0aca;
    FD1P3IX alu_b_i0_i7 (.D(float_alu_b[7]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[7]));
    defparam alu_b_i0_i7.GSR = "DISABLED";
    LUT4 mux_4232_i23_3_lut (.A(add_c[22]), .B(sub_c[22]), .C(n1148[2]), 
         .Z(n13267[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i23_3_lut.init = 16'hcaca;
    PFUMX mux_4242_i31 (.BLUT(n13267[30]), .ALUT(n13369[30]), .C0(n67175), 
          .Z(n13437[30]));
    PFUMX mux_4242_i30 (.BLUT(n13267[29]), .ALUT(n13369[29]), .C0(n67175), 
          .Z(n13437[29]));
    FD1P3IX alu_b_i0_i8 (.D(float_alu_b[8]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[8]));
    defparam alu_b_i0_i8.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(float_alu_ready), .B(n70866), .C(SDA_c), .D(n2050), 
         .Z(n4617)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_960 (.A(float_alu_ready), .B(n70866), .C(SDA_c), 
         .D(n2084), .Z(n15113)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_960.init = 16'h0200;
    FD1P3IX alu_b_i0_i9 (.D(float_alu_b[9]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[9]));
    defparam alu_b_i0_i9.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut_adj_961 (.A(float_alu_ready), .B(n70866), .C(SDA_c), 
         .D(n2072), .Z(n4599)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_961.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_962 (.A(\float_alu_mode[2] ), .B(n70850), .C(\float_alu_mode[1] ), 
         .D(n1155), .Z(n110)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_962.init = 16'hff04;
    LUT4 i1_2_lut_3_lut_rep_852 (.A(float_alu_ready), .B(n70866), .C(SDA_c), 
         .Z(n70822)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_rep_852.init = 16'h0202;
    FD1P3IX alu_b_i0_i10 (.D(float_alu_b[10]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[10]));
    defparam alu_b_i0_i10.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(float_alu_ready), .B(n70866), .C(n2036), .D(n2086), 
         .Z(n23655)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2220;
    PFUMX mux_4242_i29 (.BLUT(n13267[28]), .ALUT(n13369[28]), .C0(n67175), 
          .Z(n13437[28]));
    PFUMX mux_4242_i28 (.BLUT(n13267[27]), .ALUT(n13369[27]), .C0(n67175), 
          .Z(n13437[27]));
    FD1P3IX alu_b_i0_i11 (.D(float_alu_b[11]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[11]));
    defparam alu_b_i0_i11.GSR = "DISABLED";
    PFUMX mux_4242_i27 (.BLUT(n13267[26]), .ALUT(n13369[26]), .C0(n67175), 
          .Z(n13437[26]));
    PFUMX mux_4242_i26 (.BLUT(n13267[25]), .ALUT(n13369[25]), .C0(n67175), 
          .Z(n13437[25]));
    FD1P3IX alu_b_i0_i12 (.D(float_alu_b[12]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[12]));
    defparam alu_b_i0_i12.GSR = "DISABLED";
    PFUMX mux_4242_i25 (.BLUT(n13267[24]), .ALUT(n13369[24]), .C0(n67175), 
          .Z(n13437[24]));
    FD1P3IX alu_b_i0_i13 (.D(float_alu_b[13]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[13]));
    defparam alu_b_i0_i13.GSR = "DISABLED";
    PFUMX mux_4242_i24 (.BLUT(n13267[23]), .ALUT(n13369[23]), .C0(n67175), 
          .Z(n13437[23]));
    FD1P3IX alu_b_i0_i14 (.D(float_alu_b[14]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[14]));
    defparam alu_b_i0_i14.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i15 (.D(float_alu_b[15]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[15]));
    defparam alu_b_i0_i15.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i16 (.D(float_alu_b[16]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[16]));
    defparam alu_b_i0_i16.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i17 (.D(float_alu_b[17]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[17]));
    defparam alu_b_i0_i17.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i18 (.D(float_alu_b[18]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[18]));
    defparam alu_b_i0_i18.GSR = "DISABLED";
    FD1P3AX sub_ce_83 (.D(n23885), .SP(n23670), .CK(clock), .Q(sub_ce));
    defparam sub_ce_83.GSR = "DISABLED";
    FD1P3AX add_enable_80 (.D(n70841), .SP(n66613), .CK(clock), .Q(add_enable));
    defparam add_enable_80.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i19 (.D(float_alu_b[19]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[19]));
    defparam alu_b_i0_i19.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i20 (.D(float_alu_b[20]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[20]));
    defparam alu_b_i0_i20.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i21 (.D(float_alu_b[21]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[21]));
    defparam alu_b_i0_i21.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i22 (.D(float_alu_b[22]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[22]));
    defparam alu_b_i0_i22.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i23 (.D(float_alu_b[23]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[23]));
    defparam alu_b_i0_i23.GSR = "DISABLED";
    PFUMX mux_4242_i23 (.BLUT(n13267[22]), .ALUT(n13369[22]), .C0(n67175), 
          .Z(n13437[22]));
    FD1P3IX alu_b_i0_i24 (.D(float_alu_b[24]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[24]));
    defparam alu_b_i0_i24.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i25 (.D(float_alu_b[25]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[25]));
    defparam alu_b_i0_i25.GSR = "DISABLED";
    PFUMX mux_4242_i22 (.BLUT(n13267[21]), .ALUT(n13369[21]), .C0(n67175), 
          .Z(n13437[21]));
    PFUMX mux_4242_i21 (.BLUT(n13267[20]), .ALUT(n13369[20]), .C0(n67175), 
          .Z(n13437[20]));
    PFUMX mux_4242_i20 (.BLUT(n13267[19]), .ALUT(n13369[19]), .C0(n67175), 
          .Z(n13437[19]));
    PFUMX mux_4242_i19 (.BLUT(n13267[18]), .ALUT(n13369[18]), .C0(n67175), 
          .Z(n13437[18]));
    PFUMX mux_4242_i18 (.BLUT(n13267[17]), .ALUT(n13369[17]), .C0(n67175), 
          .Z(n13437[17]));
    LUT4 i12196_1_lut (.A(n1148[2]), .Z(n23885)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12196_1_lut.init = 16'h5555;
    FD1P3IX alu_b_i0_i26 (.D(float_alu_b[26]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[26]));
    defparam alu_b_i0_i26.GSR = "DISABLED";
    PFUMX mux_4242_i17 (.BLUT(n13267[16]), .ALUT(n13369[16]), .C0(n67175), 
          .Z(n13437[16]));
    PFUMX mux_4242_i16 (.BLUT(n13267[15]), .ALUT(n13369[15]), .C0(n67175), 
          .Z(n13437[15]));
    PFUMX mux_4242_i15 (.BLUT(n13267[14]), .ALUT(n13369[14]), .C0(n67175), 
          .Z(n13437[14]));
    PFUMX mux_4242_i14 (.BLUT(n13267[13]), .ALUT(n13369[13]), .C0(n67175), 
          .Z(n13437[13]));
    PFUMX mux_4242_i13 (.BLUT(n13267[12]), .ALUT(n13369[12]), .C0(n67175), 
          .Z(n13437[12]));
    PFUMX mux_4242_i12 (.BLUT(n13267[11]), .ALUT(n13369[11]), .C0(n67175), 
          .Z(n13437[11]));
    PFUMX mux_4242_i11 (.BLUT(n13267[10]), .ALUT(n13369[10]), .C0(n67175), 
          .Z(n13437[10]));
    PFUMX mux_4242_i10 (.BLUT(n13267[9]), .ALUT(n13369[9]), .C0(n67175), 
          .Z(n13437[9]));
    FD1P3AX alu_c_i0_i30 (.D(n13437[30]), .SP(n70744), .CK(clock), .Q(float_alu_c[30]));
    defparam alu_c_i0_i30.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i29 (.D(n13437[29]), .SP(n70744), .CK(clock), .Q(float_alu_c[29]));
    defparam alu_c_i0_i29.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i28 (.D(n13437[28]), .SP(n70744), .CK(clock), .Q(float_alu_c[28]));
    defparam alu_c_i0_i28.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i27 (.D(n13437[27]), .SP(n70744), .CK(clock), .Q(float_alu_c[27]));
    defparam alu_c_i0_i27.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i26 (.D(n13437[26]), .SP(n70744), .CK(clock), .Q(float_alu_c[26]));
    defparam alu_c_i0_i26.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i25 (.D(n13437[25]), .SP(n70744), .CK(clock), .Q(float_alu_c[25]));
    defparam alu_c_i0_i25.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i24 (.D(n13437[24]), .SP(n70744), .CK(clock), .Q(float_alu_c[24]));
    defparam alu_c_i0_i24.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i23 (.D(n13437[23]), .SP(n70744), .CK(clock), .Q(float_alu_c[23]));
    defparam alu_c_i0_i23.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i22 (.D(n13437[22]), .SP(n70744), .CK(clock), .Q(float_alu_c[22]));
    defparam alu_c_i0_i22.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i21 (.D(n13437[21]), .SP(n70744), .CK(clock), .Q(float_alu_c[21]));
    defparam alu_c_i0_i21.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i20 (.D(n13437[20]), .SP(n70744), .CK(clock), .Q(float_alu_c[20]));
    defparam alu_c_i0_i20.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i19 (.D(n13437[19]), .SP(n70744), .CK(clock), .Q(float_alu_c[19]));
    defparam alu_c_i0_i19.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i18 (.D(n13437[18]), .SP(n70744), .CK(clock), .Q(float_alu_c[18]));
    defparam alu_c_i0_i18.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i17 (.D(n13437[17]), .SP(n70744), .CK(clock), .Q(float_alu_c[17]));
    defparam alu_c_i0_i17.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i16 (.D(n13437[16]), .SP(n70744), .CK(clock), .Q(float_alu_c[16]));
    defparam alu_c_i0_i16.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i15 (.D(n13437[15]), .SP(n70744), .CK(clock), .Q(float_alu_c[15]));
    defparam alu_c_i0_i15.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i14 (.D(n13437[14]), .SP(n70744), .CK(clock), .Q(float_alu_c[14]));
    defparam alu_c_i0_i14.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i13 (.D(n13437[13]), .SP(n70744), .CK(clock), .Q(float_alu_c[13]));
    defparam alu_c_i0_i13.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i12 (.D(n13437[12]), .SP(n70744), .CK(clock), .Q(float_alu_c[12]));
    defparam alu_c_i0_i12.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i11 (.D(n13437[11]), .SP(n70744), .CK(clock), .Q(float_alu_c[11]));
    defparam alu_c_i0_i11.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i10 (.D(n13437[10]), .SP(n70744), .CK(clock), .Q(float_alu_c[10]));
    defparam alu_c_i0_i10.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i9 (.D(n13437[9]), .SP(n70744), .CK(clock), .Q(float_alu_c[9]));
    defparam alu_c_i0_i9.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i8 (.D(n13437[8]), .SP(n70744), .CK(clock), .Q(float_alu_c[8]));
    defparam alu_c_i0_i8.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i7 (.D(n13437[7]), .SP(n70744), .CK(clock), .Q(float_alu_c[7]));
    defparam alu_c_i0_i7.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i6 (.D(n13437[6]), .SP(n70744), .CK(clock), .Q(float_alu_c[6]));
    defparam alu_c_i0_i6.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i5 (.D(n13437[5]), .SP(n70744), .CK(clock), .Q(float_alu_c[5]));
    defparam alu_c_i0_i5.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i4 (.D(n13437[4]), .SP(n70744), .CK(clock), .Q(float_alu_c[4]));
    defparam alu_c_i0_i4.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i3 (.D(n13437[3]), .SP(n70744), .CK(clock), .Q(float_alu_c[3]));
    defparam alu_c_i0_i3.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i2 (.D(n13437[2]), .SP(n70744), .CK(clock), .Q(float_alu_c[2]));
    defparam alu_c_i0_i2.GSR = "DISABLED";
    FD1P3AX alu_c_i0_i1 (.D(n13437[1]), .SP(n70744), .CK(clock), .Q(float_alu_c[1]));
    defparam alu_c_i0_i1.GSR = "DISABLED";
    PFUMX mux_4242_i9 (.BLUT(n13267[8]), .ALUT(n13369[8]), .C0(n67175), 
          .Z(n13437[8]));
    PFUMX mux_4242_i8 (.BLUT(n13267[7]), .ALUT(n13369[7]), .C0(n67175), 
          .Z(n13437[7]));
    PFUMX mux_4242_i7 (.BLUT(n13267[6]), .ALUT(n13369[6]), .C0(n67175), 
          .Z(n13437[6]));
    PFUMX mux_4242_i6 (.BLUT(n13267[5]), .ALUT(n13369[5]), .C0(n67175), 
          .Z(n13437[5]));
    FD1P3IX alu_b_i0_i27 (.D(float_alu_b[27]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_b[27]));
    defparam alu_b_i0_i27.GSR = "DISABLED";
    PFUMX mux_4242_i5 (.BLUT(n13267[4]), .ALUT(n13369[4]), .C0(n67175), 
          .Z(n13437[4]));
    FD1P3IX alu_b_i0_i28 (.D(float_alu_b[28]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[28]));
    defparam alu_b_i0_i28.GSR = "DISABLED";
    PFUMX mux_4242_i4 (.BLUT(n13267[3]), .ALUT(n13369[3]), .C0(n67175), 
          .Z(n13437[3]));
    PFUMX mux_4242_i3 (.BLUT(n13267[2]), .ALUT(n13369[2]), .C0(n67175), 
          .Z(n13437[2]));
    FD1P3IX alu_b_i0_i29 (.D(float_alu_b[29]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[29]));
    defparam alu_b_i0_i29.GSR = "DISABLED";
    PFUMX mux_4242_i2 (.BLUT(n13267[1]), .ALUT(n13369[1]), .C0(n67175), 
          .Z(n13437[1]));
    FD1P3IX alu_a_i0_i31 (.D(float_alu_a[31]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[31]));
    defparam alu_a_i0_i31.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i30 (.D(float_alu_a[30]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[30]));
    defparam alu_a_i0_i30.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i29 (.D(float_alu_a[29]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[29]));
    defparam alu_a_i0_i29.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i30 (.D(float_alu_b[30]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[30]));
    defparam alu_b_i0_i30.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i28 (.D(float_alu_a[28]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[28]));
    defparam alu_a_i0_i28.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i31 (.D(float_alu_b[31]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[31]));
    defparam alu_b_i0_i31.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i27 (.D(float_alu_a[27]), .SP(n23632), .CD(n23974), 
            .CK(clock), .Q(alu_a[27]));
    defparam alu_a_i0_i27.GSR = "DISABLED";
    LUT4 mux_4234_i24_3_lut (.A(mul_c[23]), .B(div_c[23]), .C(n1148[4]), 
         .Z(n13301[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i24_3_lut.init = 16'hcaca;
    LUT4 i54851_4_lut (.A(n13301[23]), .B(eR_e3[0]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[23])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54851_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i24_3_lut (.A(add_c[23]), .B(sub_c[23]), .C(n1148[2]), 
         .Z(n13267[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i24_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i25_3_lut (.A(mul_c[24]), .B(div_c[24]), .C(n1148[4]), 
         .Z(n13301[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i25_3_lut.init = 16'hcaca;
    FD1P3IX alu_a_i0_i26 (.D(float_alu_a[26]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[26]));
    defparam alu_a_i0_i26.GSR = "DISABLED";
    LUT4 i54849_4_lut (.A(n13301[24]), .B(eR_e3[1]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[24])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54849_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i25_3_lut (.A(add_c[24]), .B(sub_c[24]), .C(n1148[2]), 
         .Z(n13267[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i25_3_lut.init = 16'hcaca;
    FD1P3IX alu_a_i0_i25 (.D(float_alu_a[25]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[25]));
    defparam alu_a_i0_i25.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i24 (.D(float_alu_a[24]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[24]));
    defparam alu_a_i0_i24.GSR = "DISABLED";
    PFUMX mux_4242_i1 (.BLUT(n13267[0]), .ALUT(n13369[0]), .C0(n67175), 
          .Z(n13437[0]));
    FD1P3IX alu_a_i0_i23 (.D(float_alu_a[23]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[23]));
    defparam alu_a_i0_i23.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i22 (.D(float_alu_a[22]), .SP(n23632), .CD(n23974), 
            .CK(clock), .Q(alu_a[22]));
    defparam alu_a_i0_i22.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i21 (.D(float_alu_a[21]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[21]));
    defparam alu_a_i0_i21.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i20 (.D(float_alu_a[20]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[20]));
    defparam alu_a_i0_i20.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i19 (.D(float_alu_a[19]), .SP(n23632), .CD(n23974), 
            .CK(clock), .Q(alu_a[19]));
    defparam alu_a_i0_i19.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i18 (.D(float_alu_a[18]), .SP(n23632), .CD(n73820), 
            .CK(clock), .Q(alu_a[18]));
    defparam alu_a_i0_i18.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i17 (.D(float_alu_a[17]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[17]));
    defparam alu_a_i0_i17.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i16 (.D(float_alu_a[16]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[16]));
    defparam alu_a_i0_i16.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i15 (.D(float_alu_a[15]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[15]));
    defparam alu_a_i0_i15.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i14 (.D(float_alu_a[14]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_a[14]));
    defparam alu_a_i0_i14.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i13 (.D(float_alu_a[13]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[13]));
    defparam alu_a_i0_i13.GSR = "DISABLED";
    LUT4 mux_4234_i26_3_lut (.A(mul_c[25]), .B(div_c[25]), .C(n1148[4]), 
         .Z(n13301[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i26_3_lut.init = 16'hcaca;
    LUT4 i54847_4_lut (.A(n13301[25]), .B(eR_e3[2]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[25])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54847_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i26_3_lut (.A(add_c[25]), .B(sub_c[25]), .C(n1148[2]), 
         .Z(n13267[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i26_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i27_3_lut (.A(mul_c[26]), .B(div_c[26]), .C(n1148[4]), 
         .Z(n13301[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i27_3_lut.init = 16'hcaca;
    LUT4 i54845_4_lut (.A(n13301[26]), .B(eR_e3[3]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[26])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54845_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i27_3_lut (.A(add_c[26]), .B(sub_c[26]), .C(n1148[2]), 
         .Z(n13267[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i27_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i28_3_lut (.A(mul_c[27]), .B(div_c[27]), .C(n1148[4]), 
         .Z(n13301[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i28_3_lut.init = 16'hcaca;
    LUT4 i54843_4_lut (.A(n13301[27]), .B(eR_e3[4]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[27])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54843_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i28_3_lut (.A(add_c[27]), .B(sub_c[27]), .C(n1148[2]), 
         .Z(n13267[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i28_3_lut.init = 16'hcaca;
    FD1P3IX alu_c_i0_i31 (.D(n13369[31]), .SP(n70744), .CD(n23979), .CK(clock), 
            .Q(float_alu_c[31]));
    defparam alu_c_i0_i31.GSR = "DISABLED";
    LUT4 i1_2_lut_2_lut_3_lut (.A(n70866), .B(n1156), .C(n73809), .Z(n45611)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'h8f8f;
    LUT4 mux_4234_i29_3_lut (.A(mul_c[28]), .B(div_c[28]), .C(n1148[4]), 
         .Z(n13301[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i29_3_lut.init = 16'hcaca;
    LUT4 i54841_4_lut (.A(n13301[28]), .B(eR_e3[5]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[28])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54841_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i29_3_lut (.A(add_c[28]), .B(sub_c[28]), .C(n1148[2]), 
         .Z(n13267[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i29_3_lut.init = 16'hcaca;
    LUT4 i55044_4_lut_rep_808 (.A(wait_counter[17]), .B(n14), .C(n10), 
         .D(wait_counter[21]), .Z(n70778)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i55044_4_lut_rep_808.init = 16'h0001;
    LUT4 i1_3_lut_4_lut_adj_963 (.A(n73809), .B(SDA_c), .C(n70814), .D(n1148[4]), 
         .Z(n142_adj_528)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_963.init = 16'h2220;
    LUT4 i1_3_lut_4_lut_adj_964 (.A(n73809), .B(SDA_c), .C(n1148[3]), 
         .D(n70790), .Z(n141)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_964.init = 16'h2220;
    LUT4 i1_3_lut_4_lut_adj_965 (.A(n73809), .B(SDA_c), .C(n1148[2]), 
         .D(n70781), .Z(n23670)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_965.init = 16'h2220;
    LUT4 i177_2_lut_rep_797 (.A(n73809), .B(SDA_c), .Z(n70767)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i177_2_lut_rep_797.init = 16'hdddd;
    LUT4 i23551_4_lut (.A(n70788), .B(n130[30]), .C(n73809), .D(wait_counter[30]), 
         .Z(n23850)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23551_4_lut.init = 16'hac0c;
    LUT4 i23548_4_lut (.A(n70788), .B(n130[29]), .C(n73809), .D(wait_counter[29]), 
         .Z(n23854)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23548_4_lut.init = 16'hac0c;
    LUT4 i23557_4_lut (.A(n70788), .B(n130[28]), .C(n73809), .D(wait_counter[28]), 
         .Z(n23856)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23557_4_lut.init = 16'hac0c;
    LUT4 i23560_4_lut (.A(n70788), .B(n130[27]), .C(n73809), .D(wait_counter[27]), 
         .Z(n23858)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23560_4_lut.init = 16'hac0c;
    LUT4 i23554_4_lut (.A(n70788), .B(n130[26]), .C(n73809), .D(wait_counter[26]), 
         .Z(n23860)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23554_4_lut.init = 16'hac0c;
    LUT4 i12173_4_lut (.A(n70788), .B(n130[25]), .C(n73809), .D(wait_counter[25]), 
         .Z(n23862)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12173_4_lut.init = 16'hac0c;
    LUT4 i23491_4_lut (.A(n70788), .B(n130[24]), .C(n73809), .D(wait_counter[24]), 
         .Z(n23871)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23491_4_lut.init = 16'hac0c;
    LUT4 i23488_4_lut (.A(n70788), .B(n130[23]), .C(n73809), .D(wait_counter[23]), 
         .Z(n23877)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23488_4_lut.init = 16'hac0c;
    LUT4 i23494_4_lut (.A(n70788), .B(n130[22]), .C(n73809), .D(wait_counter[22]), 
         .Z(n23882)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23494_4_lut.init = 16'hac0c;
    LUT4 i23485_4_lut (.A(n70788), .B(n130[21]), .C(n73809), .D(wait_counter[21]), 
         .Z(n23884)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23485_4_lut.init = 16'hac0c;
    LUT4 i23475_4_lut (.A(n70788), .B(n130[20]), .C(n73809), .D(wait_counter[20]), 
         .Z(n23891)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23475_4_lut.init = 16'hac0c;
    LUT4 i12204_4_lut (.A(n70788), .B(n130[19]), .C(n73809), .D(wait_counter[19]), 
         .Z(n23893)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12204_4_lut.init = 16'hac0c;
    LUT4 i12206_4_lut (.A(n70788), .B(n130[18]), .C(n73809), .D(wait_counter[18]), 
         .Z(n23895)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12206_4_lut.init = 16'hac0c;
    LUT4 i23500_4_lut (.A(n70788), .B(n130[17]), .C(n73809), .D(wait_counter[17]), 
         .Z(n23897)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i23500_4_lut.init = 16'hac0c;
    LUT4 i12210_4_lut (.A(n70788), .B(n130[16]), .C(n73809), .D(wait_counter[16]), 
         .Z(n23899)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12210_4_lut.init = 16'hac0c;
    LUT4 i12212_4_lut (.A(n70788), .B(n130[15]), .C(n73809), .D(wait_counter[15]), 
         .Z(n23901)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12212_4_lut.init = 16'hac0c;
    LUT4 i12214_4_lut (.A(n70788), .B(n130[14]), .C(n73809), .D(wait_counter[14]), 
         .Z(n23903)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12214_4_lut.init = 16'hac0c;
    LUT4 i33877_4_lut (.A(n70788), .B(n130[13]), .C(n73809), .D(wait_counter[13]), 
         .Z(n23905)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i33877_4_lut.init = 16'hac0c;
    LUT4 i33875_4_lut (.A(n70788), .B(n130[12]), .C(n73809), .D(wait_counter[12]), 
         .Z(n23911)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i33875_4_lut.init = 16'hac0c;
    LUT4 i12224_4_lut (.A(n70788), .B(n130[11]), .C(n73809), .D(wait_counter[11]), 
         .Z(n23913)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12224_4_lut.init = 16'hac0c;
    LUT4 i12178_4_lut (.A(n70788), .B(n130[10]), .C(n73809), .D(wait_counter[10]), 
         .Z(n23867)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12178_4_lut.init = 16'hac0c;
    LUT4 i12184_4_lut (.A(n70788), .B(n130[9]), .C(n73809), .D(wait_counter[9]), 
         .Z(n23873)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12184_4_lut.init = 16'hac0c;
    LUT4 i12228_4_lut (.A(n70788), .B(n130[6]), .C(n73809), .D(wait_counter[6]), 
         .Z(n23917)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12228_4_lut.init = 16'hac0c;
    LUT4 i12230_4_lut (.A(n70788), .B(n130[5]), .C(n73809), .D(wait_counter[5]), 
         .Z(n23919)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12230_4_lut.init = 16'hac0c;
    LUT4 i12232_4_lut (.A(n70788), .B(n130[4]), .C(n73809), .D(wait_counter[4]), 
         .Z(n23921)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i12232_4_lut.init = 16'hac0c;
    LUT4 i53905_2_lut (.A(\float_alu_mode[2] ), .B(float_alu_mode[0]), .Z(n66808)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53905_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(\float_alu_mode[1] ), .B(n130[1]), .C(n73809), 
         .D(n66808), .Z(n65745)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A !(B+(C)))) */ ;
    defparam i22_4_lut.init = 16'h5cfc;
    LUT4 mux_4234_i30_3_lut (.A(mul_c[29]), .B(div_c[29]), .C(n1148[4]), 
         .Z(n13301[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i30_3_lut.init = 16'hcaca;
    LUT4 i54839_4_lut (.A(n13301[29]), .B(eR_e3[6]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[29])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i54839_4_lut.init = 16'hfaca;
    LUT4 mux_4232_i30_3_lut (.A(add_c[29]), .B(sub_c[29]), .C(n1148[2]), 
         .Z(n13267[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i30_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n73818), .B(n2086), .C(n2036), .D(n2082), .Z(n23653)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'haaa8;
    LUT4 mux_4234_i31_3_lut (.A(mul_c[30]), .B(div_c[30]), .C(n1148[4]), 
         .Z(n13301[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i31_3_lut.init = 16'hcaca;
    LUT4 i54837_4_lut (.A(n13301[30]), .B(eR_e3[7]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54837_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i31_3_lut (.A(add_c[30]), .B(sub_c[30]), .C(n1148[2]), 
         .Z(n13267[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i31_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(n73809), .B(n1156), .C(n142), .D(SDA_c), 
         .Z(n66613)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 i37_3_lut_3_lut (.A(n73809), .B(n130[3]), .C(n47), .Z(n163[3])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i37_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_2_lut (.A(n73809), .B(n130[7]), .Z(n23915)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_966 (.A(n73809), .B(n130[8]), .Z(n23875)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_2_lut_adj_966.init = 16'h4444;
    LUT4 i1_4_lut_adj_967 (.A(SDA_c), .B(n73809), .C(n45598), .D(n110), 
         .Z(n23819)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_967.init = 16'h5450;
    FD1P3IX alu_a_i0_i12 (.D(float_alu_a[12]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[12]));
    defparam alu_a_i0_i12.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i31 (.D(n63068), .SP(n70716), .CK(clock), .Q(float_alu_a[31]));
    defparam float_alu_a_i0_i31.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i30 (.D(n62958), .SP(n70716), .CK(clock), .Q(float_alu_a[30]));
    defparam float_alu_a_i0_i30.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i27 (.D(n66522), .SP(n70716), .CK(clock), .Q(float_alu_a[27]));
    defparam float_alu_a_i0_i27.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i25 (.D(n66524), .SP(n70716), .CK(clock), .Q(float_alu_a[25]));
    defparam float_alu_a_i0_i25.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i23 (.D(n63156), .SP(n70716), .CK(clock), .Q(float_alu_a[23]));
    defparam float_alu_a_i0_i23.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i22 (.D(n63069), .SP(n70716), .CK(clock), .Q(float_alu_a[22]));
    defparam float_alu_a_i0_i22.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i21 (.D(n63070), .SP(n70716), .CK(clock), .Q(float_alu_a[21]));
    defparam float_alu_a_i0_i21.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i20 (.D(n62961), .SP(n70716), .CK(clock), .Q(float_alu_a[20]));
    defparam float_alu_a_i0_i20.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i19 (.D(n63102), .SP(n70716), .CK(clock), .Q(float_alu_a[19]));
    defparam float_alu_a_i0_i19.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i18 (.D(n63103), .SP(n70716), .CK(clock), .Q(float_alu_a[18]));
    defparam float_alu_a_i0_i18.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i17 (.D(n63104), .SP(n70716), .CK(clock), .Q(float_alu_a[17]));
    defparam float_alu_a_i0_i17.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i16 (.D(n63106), .SP(n70716), .CK(clock), .Q(float_alu_a[16]));
    defparam float_alu_a_i0_i16.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i15 (.D(n63105), .SP(n70716), .CK(clock), .Q(float_alu_a[15]));
    defparam float_alu_a_i0_i15.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i14 (.D(n63107), .SP(n70716), .CK(clock), .Q(float_alu_a[14]));
    defparam float_alu_a_i0_i14.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i13 (.D(n63114), .SP(n70716), .CK(clock), .Q(float_alu_a[13]));
    defparam float_alu_a_i0_i13.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i12 (.D(n63109), .SP(n70716), .CK(clock), .Q(float_alu_a[12]));
    defparam float_alu_a_i0_i12.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i11 (.D(n63115), .SP(n70716), .CK(clock), .Q(float_alu_a[11]));
    defparam float_alu_a_i0_i11.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i10 (.D(n63116), .SP(n70716), .CK(clock), .Q(float_alu_a[10]));
    defparam float_alu_a_i0_i10.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i9 (.D(n63120), .SP(n70716), .CK(clock), .Q(float_alu_a[9]));
    defparam float_alu_a_i0_i9.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i8 (.D(n63122), .SP(n70716), .CK(clock), .Q(float_alu_a[8]));
    defparam float_alu_a_i0_i8.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i7 (.D(n63128), .SP(n70716), .CK(clock), .Q(float_alu_a[7]));
    defparam float_alu_a_i0_i7.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i6 (.D(n63131), .SP(n70716), .CK(clock), .Q(float_alu_a[6]));
    defparam float_alu_a_i0_i6.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i5 (.D(n63139), .SP(n70716), .CK(clock), .Q(float_alu_a[5]));
    defparam float_alu_a_i0_i5.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i4 (.D(n63147), .SP(n70716), .CK(clock), .Q(float_alu_a[4]));
    defparam float_alu_a_i0_i4.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i3 (.D(n63150), .SP(n70716), .CK(clock), .Q(float_alu_a[3]));
    defparam float_alu_a_i0_i3.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i2 (.D(n62964), .SP(n70716), .CK(clock), .Q(float_alu_a[2]));
    defparam float_alu_a_i0_i2.GSR = "DISABLED";
    FD1P3AX float_alu_a_i0_i1 (.D(n62966), .SP(n70716), .CK(clock), .Q(float_alu_a[1]));
    defparam float_alu_a_i0_i1.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i11 (.D(float_alu_a[11]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_a[11]));
    defparam alu_a_i0_i11.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i10 (.D(float_alu_a[10]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[10]));
    defparam alu_a_i0_i10.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i9 (.D(float_alu_a[9]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[9]));
    defparam alu_a_i0_i9.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i8 (.D(float_alu_a[8]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[8]));
    defparam alu_a_i0_i8.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i7 (.D(float_alu_a[7]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[7]));
    defparam alu_a_i0_i7.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i6 (.D(float_alu_a[6]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_a[6]));
    defparam alu_a_i0_i6.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i5 (.D(float_alu_a[5]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[5]));
    defparam alu_a_i0_i5.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i4 (.D(float_alu_a[4]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[4]));
    defparam alu_a_i0_i4.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i3 (.D(float_alu_a[3]), .SP(n73817), .CD(n23974), 
            .CK(clock), .Q(alu_a[3]));
    defparam alu_a_i0_i3.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i2 (.D(float_alu_a[2]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[2]));
    defparam alu_a_i0_i2.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i1 (.D(float_alu_a[1]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[1]));
    defparam alu_a_i0_i1.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i31 (.D(float_alu_a[31]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(mXs_0[24]));
    defparam exp_a_i0_i31.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i30 (.D(float_alu_a[30]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[30]));
    defparam exp_a_i0_i30.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i29 (.D(float_alu_a[29]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[29]));
    defparam exp_a_i0_i29.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i28 (.D(float_alu_a[28]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[28]));
    defparam exp_a_i0_i28.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i27 (.D(float_alu_a[27]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[27]));
    defparam exp_a_i0_i27.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i26 (.D(float_alu_a[26]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[26]));
    defparam exp_a_i0_i26.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i25 (.D(float_alu_a[25]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[25]));
    defparam exp_a_i0_i25.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i24 (.D(float_alu_a[24]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[24]));
    defparam exp_a_i0_i24.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i23 (.D(float_alu_a[23]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[23]));
    defparam exp_a_i0_i23.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i22 (.D(float_alu_a[22]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[22]));
    defparam exp_a_i0_i22.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i21 (.D(float_alu_a[21]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[21]));
    defparam exp_a_i0_i21.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i20 (.D(float_alu_a[20]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[20]));
    defparam exp_a_i0_i20.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i19 (.D(float_alu_a[19]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[19]));
    defparam exp_a_i0_i19.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i18 (.D(float_alu_a[18]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[18]));
    defparam exp_a_i0_i18.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i17 (.D(float_alu_a[17]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[17]));
    defparam exp_a_i0_i17.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i16 (.D(float_alu_a[16]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[16]));
    defparam exp_a_i0_i16.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i15 (.D(float_alu_a[15]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[15]));
    defparam exp_a_i0_i15.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i14 (.D(float_alu_a[14]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[14]));
    defparam exp_a_i0_i14.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i13 (.D(float_alu_a[13]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[13]));
    defparam exp_a_i0_i13.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i12 (.D(float_alu_a[12]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[12]));
    defparam exp_a_i0_i12.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i11 (.D(float_alu_a[11]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[11]));
    defparam exp_a_i0_i11.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i10 (.D(float_alu_a[10]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[10]));
    defparam exp_a_i0_i10.GSR = "DISABLED";
    FD1P3DX state_FSM__i6 (.D(n66655), .SP(n70778), .CK(clock), .CD(SDA_c), 
            .Q(n1151));
    defparam state_FSM__i6.GSR = "DISABLED";
    FD1P3DX state_FSM__i5 (.D(n22189), .SP(n70778), .CK(clock), .CD(SDA_c), 
            .Q(n1148[4]));
    defparam state_FSM__i5.GSR = "DISABLED";
    FD1P3DX state_FSM__i4 (.D(n22185), .SP(n70778), .CK(clock), .CD(SDA_c), 
            .Q(n1148[3]));
    defparam state_FSM__i4.GSR = "DISABLED";
    FD1P3DX state_FSM__i3 (.D(n22187), .SP(n70778), .CK(clock), .CD(SDA_c), 
            .Q(n1148[2]));
    defparam state_FSM__i3.GSR = "DISABLED";
    FD1P3DX state_FSM__i2 (.D(n70793), .SP(n70778), .CK(clock), .CD(SDA_c), 
            .Q(n1155));
    defparam state_FSM__i2.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i9 (.D(float_alu_a[9]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[9]));
    defparam exp_a_i0_i9.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i8 (.D(float_alu_a[8]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[8]));
    defparam exp_a_i0_i8.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i7 (.D(float_alu_a[7]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[7]));
    defparam exp_a_i0_i7.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i6 (.D(float_alu_a[6]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[6]));
    defparam exp_a_i0_i6.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i5 (.D(float_alu_a[5]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[5]));
    defparam exp_a_i0_i5.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i4 (.D(float_alu_a[4]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[4]));
    defparam exp_a_i0_i4.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i3 (.D(float_alu_a[3]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[3]));
    defparam exp_a_i0_i3.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i2 (.D(float_alu_a[2]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[2]));
    defparam exp_a_i0_i2.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i1 (.D(float_alu_a[1]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[1]));
    defparam exp_a_i0_i1.GSR = "DISABLED";
    LUT4 i2_1_lut (.A(\float_alu_mode[1] ), .Z(n45720)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut.init = 16'h5555;
    LUT4 i1_2_lut (.A(SDA_c), .B(n1673), .Z(n4445)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i6_4_lut_adj_968 (.A(wait_counter[5]), .B(wait_counter[29]), .C(wait_counter[7]), 
         .D(wait_counter[8]), .Z(n16_adj_531)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_968.init = 16'hfffe;
    LUT4 i7_4_lut (.A(wait_counter[28]), .B(wait_counter[26]), .C(wait_counter[27]), 
         .D(wait_counter[30]), .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i9_4_lut_adj_969 (.A(n17), .B(wait_counter[1]), .C(n16_adj_531), 
         .D(wait_counter[0]), .Z(n66700)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_adj_969.init = 16'hfffe;
    LUT4 i5_2_lut (.A(wait_counter[11]), .B(wait_counter[15]), .Z(n20)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(wait_counter[2]), .B(wait_counter[19]), .C(wait_counter[3]), 
         .D(wait_counter[12]), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_970 (.A(wait_counter[16]), .B(wait_counter[10]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_970.init = 16'heeee;
    FD1P3AX exp_a_i0_i32 (.D(n45720), .SP(n23722), .CK(clock), .Q(exp_a[32]));
    defparam exp_a_i0_i32.GSR = "DISABLED";
    LUT4 i5_4_lut (.A(n139_adj_532), .B(wait_counter[17]), .C(wait_counter[24]), 
         .D(wait_counter[23]), .Z(n12)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i5_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_adj_971 (.A(SDA_c), .B(n1156), .Z(n4_c)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_971.init = 16'h4444;
    LUT4 i6_4_lut_adj_972 (.A(wait_counter[22]), .B(n12), .C(wait_counter[20]), 
         .D(wait_counter[21]), .Z(n66575)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i6_4_lut_adj_972.init = 16'h0004;
    LUT4 i12284_4_lut (.A(n73816), .B(n66208), .C(n66575), .D(n4_c), 
         .Z(n23974)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;
    defparam i12284_4_lut.init = 16'h8aaa;
    FD1P3DX wait_counter_4646_4647__i1 (.D(n69007), .SP(n45611), .CK(clock), 
            .CD(SDA_c), .Q(wait_counter[0]));
    defparam wait_counter_4646_4647__i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(\float_alu_mode[1] ), .B(n70767), .C(n70856), .D(n1156), 
         .Z(n23632)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;
    defparam i2_4_lut.init = 16'h3200;
    FD1P3DX wait_counter_4646_4647__i2 (.D(n65745), .SP(n45611), .CK(clock), 
            .CD(SDA_c), .Q(wait_counter[1]));
    defparam wait_counter_4646_4647__i2.GSR = "DISABLED";
    FD1P3AX mul_ce_85 (.D(n1442), .SP(n141), .CK(clock), .Q(mul_ce));
    defparam mul_ce_85.GSR = "DISABLED";
    FD1P3DX float_alu_mode_i0_i0 (.D(n23942), .SP(n27939), .CK(clock), 
            .CD(SDA_c), .Q(float_alu_mode[0]));
    defparam float_alu_mode_i0_i0.GSR = "DISABLED";
    FD1P3IX alu_b_i0_i0 (.D(float_alu_b[0]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_b[0]));
    defparam alu_b_i0_i0.GSR = "DISABLED";
    FD1P3DX wait_counter_4646_4647__i3 (.D(n68796), .SP(n45611), .CK(clock), 
            .CD(SDA_c), .Q(wait_counter[2]));
    defparam wait_counter_4646_4647__i3.GSR = "DISABLED";
    FD1P3DX wait_counter_4646_4647__i4 (.D(n163[3]), .SP(n45611), .CK(clock), 
            .CD(SDA_c), .Q(wait_counter[3]));
    defparam wait_counter_4646_4647__i4.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i5 (.D(n23921), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[4]));
    defparam wait_counter_4646_4647__i5.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i6 (.D(n23919), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[5]));
    defparam wait_counter_4646_4647__i6.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i7 (.D(n23917), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[6]));
    defparam wait_counter_4646_4647__i7.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i8 (.D(n23915), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[7]));
    defparam wait_counter_4646_4647__i8.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i9 (.D(n23875), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[8]));
    defparam wait_counter_4646_4647__i9.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i10 (.D(n23873), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[9]));
    defparam wait_counter_4646_4647__i10.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i11 (.D(n23867), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[10]));
    defparam wait_counter_4646_4647__i11.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i12 (.D(n23913), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[11]));
    defparam wait_counter_4646_4647__i12.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i13 (.D(n23911), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[12]));
    defparam wait_counter_4646_4647__i13.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i14 (.D(n23905), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[13]));
    defparam wait_counter_4646_4647__i14.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i15 (.D(n23903), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[14]));
    defparam wait_counter_4646_4647__i15.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i16 (.D(n23901), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[15]));
    defparam wait_counter_4646_4647__i16.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i17 (.D(n23899), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[16]));
    defparam wait_counter_4646_4647__i17.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i18 (.D(n23897), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[17]));
    defparam wait_counter_4646_4647__i18.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i19 (.D(n23895), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[18]));
    defparam wait_counter_4646_4647__i19.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i20 (.D(n23893), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[19]));
    defparam wait_counter_4646_4647__i20.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i21 (.D(n23891), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[20]));
    defparam wait_counter_4646_4647__i21.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i22 (.D(n23884), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[21]));
    defparam wait_counter_4646_4647__i22.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i23 (.D(n23882), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[22]));
    defparam wait_counter_4646_4647__i23.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i24 (.D(n23877), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[23]));
    defparam wait_counter_4646_4647__i24.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i25 (.D(n23871), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[24]));
    defparam wait_counter_4646_4647__i25.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i26 (.D(n23862), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[25]));
    defparam wait_counter_4646_4647__i26.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i27 (.D(n23860), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[26]));
    defparam wait_counter_4646_4647__i27.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i28 (.D(n23858), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[27]));
    defparam wait_counter_4646_4647__i28.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i29 (.D(n23856), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[28]));
    defparam wait_counter_4646_4647__i29.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i30 (.D(n23854), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[29]));
    defparam wait_counter_4646_4647__i30.GSR = "DISABLED";
    FD1S3DX wait_counter_4646_4647__i31 (.D(n23850), .CK(clock), .CD(SDA_c), 
            .Q(wait_counter[30]));
    defparam wait_counter_4646_4647__i31.GSR = "DISABLED";
    FD1P3IX alu_a_i0_i0 (.D(float_alu_a[0]), .SP(n73817), .CD(n73820), 
            .CK(clock), .Q(alu_a[0]));
    defparam alu_a_i0_i0.GSR = "DISABLED";
    FD1P3AX div_ce_86 (.D(n86), .SP(n142_adj_528), .CK(clock), .Q(div_ce));
    defparam div_ce_86.GSR = "DISABLED";
    FD1P3AX add_ce_79_rep_906 (.D(n124), .SP(n23819), .CK(clock), .Q(n73804));
    defparam add_ce_79_rep_906.GSR = "DISABLED";
    FD1P3IX exp_a_i0_i0 (.D(float_alu_a[0]), .SP(n23722), .CD(n23972), 
            .CK(clock), .Q(exp_a[0]));
    defparam exp_a_i0_i0.GSR = "DISABLED";
    FD1P3JX float_alu_a_i0_i26 (.D(n63112), .SP(n70716), .PD(n24013), 
            .CK(clock), .Q(float_alu_a[26]));
    defparam float_alu_a_i0_i26.GSR = "DISABLED";
    FD1P3JX float_alu_a_i0_i24 (.D(n63111), .SP(n70716), .PD(n24013), 
            .CK(clock), .Q(float_alu_a[24]));
    defparam float_alu_a_i0_i24.GSR = "DISABLED";
    LUT4 i12282_2_lut (.A(n23722), .B(\float_alu_mode[1] ), .Z(n23972)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12282_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_973 (.A(SDA_c), .B(n73809), .C(n45598), .D(n70815), 
         .Z(n23722)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_973.init = 16'h5450;
    LUT4 mux_4234_i32_3_lut (.A(mul_c[31]), .B(div_c[31]), .C(n1148[4]), 
         .Z(n13301[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i32_3_lut.init = 16'hcaca;
    LUT4 mux_4232_i32_3_lut (.A(add_c[31]), .B(sub_c[31]), .C(n1148[2]), 
         .Z(n13267[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i32_3_lut.init = 16'hcaca;
    LUT4 i55074_2_lut_rep_846_4_lut (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .D(float_alu_ready), .Z(n70816)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i55074_2_lut_rep_846_4_lut.init = 16'h0100;
    LUT4 i55089_2_lut_rep_818_4_lut (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .D(n1156), .Z(n70788)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;
    defparam i55089_2_lut_rep_818_4_lut.init = 16'h01ff;
    FD1P3AX add_ce_79_rep_905 (.D(n124), .SP(n23819), .CK(clock), .Q(n73803));
    defparam add_ce_79_rep_905.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .D(n1156), .Z(n113)) /* synthesis lut_function=(A (B+!(D))+!A !(B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h89ff;
    LUT4 i2_3_lut_rep_896 (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .Z(n70866)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_896.init = 16'hfefe;
    LUT4 n161_bdd_3_lut (.A(n130[0]), .B(n69006), .C(n73809), .Z(n69007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n161_bdd_3_lut.init = 16'hcaca;
    LUT4 n538_bdd_3_lut (.A(\float_alu_mode[2] ), .B(float_alu_mode[0]), 
         .C(\float_alu_mode[1] ), .Z(n69006)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;
    defparam n538_bdd_3_lut.init = 16'h5c5c;
    PFUMX mux_4238_i32 (.BLUT(n13267[31]), .ALUT(n13301[31]), .C0(n70849), 
          .Z(n13369[31]));
    LUT4 i126_4_lut_4_lut (.A(float_alu_mode[0]), .B(\float_alu_mode[2] ), 
         .C(\float_alu_mode[1] ), .D(n66700), .Z(n139_adj_532)) /* synthesis lut_function=(!(A (B+(D))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i126_4_lut_4_lut.init = 16'h0036;
    LUT4 i25_2_lut_rep_886 (.A(float_alu_mode[0]), .B(\float_alu_mode[2] ), 
         .Z(n70856)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i25_2_lut_rep_886.init = 16'h6666;
    LUT4 float_alu_mode_2__bdd_3_lut (.A(\float_alu_mode[2] ), .B(float_alu_mode[0]), 
         .C(\float_alu_mode[1] ), .Z(n68795)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)))) */ ;
    defparam float_alu_mode_2__bdd_3_lut.init = 16'h1d1d;
    LUT4 n159_bdd_3_lut (.A(n130[2]), .B(n68795), .C(n73809), .Z(n68796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n159_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_974 (.A(float_alu_mode[0]), .B(n1156), 
         .C(\float_alu_mode[1] ), .D(\float_alu_mode[2] ), .Z(n66655)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_974.init = 16'h0800;
    LUT4 i1_2_lut_rep_845_3_lut (.A(float_alu_mode[0]), .B(n1156), .C(\float_alu_mode[2] ), 
         .Z(n70815)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_845_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_rep_823_4_lut (.A(float_alu_mode[0]), .B(n1156), 
         .C(\float_alu_mode[1] ), .D(\float_alu_mode[2] ), .Z(n70793)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_rep_823_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_975 (.A(float_alu_mode[0]), .B(n1156), 
         .C(\float_alu_mode[1] ), .D(\float_alu_mode[2] ), .Z(n22185)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_975.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_976 (.A(float_alu_mode[0]), .B(n1156), 
         .C(n1148[3]), .D(\float_alu_mode[1] ), .Z(n1442)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_976.init = 16'h0800;
    LUT4 i1_2_lut_rep_820_3_lut (.A(float_alu_mode[0]), .B(n1156), .C(\float_alu_mode[1] ), 
         .Z(n70790)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_820_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_880 (.A(float_alu_mode[0]), .B(n1156), .Z(n70850)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_880.init = 16'h8888;
    LUT4 i55090_2_lut_3_lut (.A(n1148[4]), .B(n1148[3]), .C(n1151), .Z(n67175)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i55090_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_879 (.A(n1148[4]), .B(n1148[3]), .Z(n70849)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_879.init = 16'heeee;
    LUT4 i12284_4_lut_rep_922 (.A(n73816), .B(n66208), .C(n66575), .D(n4_c), 
         .Z(n73820)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;
    defparam i12284_4_lut_rep_922.init = 16'h8aaa;
    CCU2D wait_counter_4646_4647_add_4_31 (.A0(wait_counter[29]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[30]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62758), .S0(n130[29]), .S1(n130[30]));
    defparam wait_counter_4646_4647_add_4_31.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_31.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_31.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_31.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_29 (.A0(wait_counter[27]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[28]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62757), .COUT(n62758), .S0(n130[27]), 
          .S1(n130[28]));
    defparam wait_counter_4646_4647_add_4_29.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_29.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_29.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_29.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_27 (.A0(wait_counter[25]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[26]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62756), .COUT(n62757), .S0(n130[25]), 
          .S1(n130[26]));
    defparam wait_counter_4646_4647_add_4_27.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_27.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_27.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_27.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_25 (.A0(wait_counter[23]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[24]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62755), .COUT(n62756), .S0(n130[23]), 
          .S1(n130[24]));
    defparam wait_counter_4646_4647_add_4_25.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_25.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_25.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_25.INJECT1_1 = "NO";
    LUT4 i55074_2_lut_rep_920 (.A(\float_alu_mode[2] ), .B(\float_alu_mode[1] ), 
         .C(float_alu_mode[0]), .D(float_alu_ready), .Z(n73818)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i55074_2_lut_rep_920.init = 16'h0100;
    LUT4 i2_4_lut_rep_919 (.A(\float_alu_mode[1] ), .B(n70767), .C(n70856), 
         .D(n1156), .Z(n73817)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;
    defparam i2_4_lut_rep_919.init = 16'h3200;
    CCU2D wait_counter_4646_4647_add_4_23 (.A0(wait_counter[21]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[22]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62754), .COUT(n62755), .S0(n130[21]), 
          .S1(n130[22]));
    defparam wait_counter_4646_4647_add_4_23.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_23.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_23.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_23.INJECT1_1 = "NO";
    LUT4 i2_4_lut_rep_918 (.A(\float_alu_mode[1] ), .B(n70767), .C(n70856), 
         .D(n1156), .Z(n73816)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;
    defparam i2_4_lut_rep_918.init = 16'h3200;
    FD1P3AX div_ce_86_rep_917 (.D(n86), .SP(n142_adj_528), .CK(clock), 
            .Q(n73815));
    defparam div_ce_86_rep_917.GSR = "DISABLED";
    CCU2D wait_counter_4646_4647_add_4_21 (.A0(wait_counter[19]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[20]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62753), .COUT(n62754), .S0(n130[19]), 
          .S1(n130[20]));
    defparam wait_counter_4646_4647_add_4_21.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_21.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_21.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_977 (.A(n73812), .B(n41808), .C(n42941), .D(n42934), 
         .Z(n25583)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_977.init = 16'ha2a0;
    CCU2D wait_counter_4646_4647_add_4_19 (.A0(wait_counter[17]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[18]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62752), .COUT(n62753), .S0(n130[17]), 
          .S1(n130[18]));
    defparam wait_counter_4646_4647_add_4_19.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_19.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_19.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_19.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_17 (.A0(wait_counter[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[16]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62751), .COUT(n62752), .S0(n130[15]), 
          .S1(n130[16]));
    defparam wait_counter_4646_4647_add_4_17.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_17.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_17.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_17.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_15 (.A0(wait_counter[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[14]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62750), .COUT(n62751), .S0(n130[13]), 
          .S1(n130[14]));
    defparam wait_counter_4646_4647_add_4_15.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_15.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_15.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_15.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_13 (.A0(wait_counter[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[12]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62749), .COUT(n62750), .S0(n130[11]), 
          .S1(n130[12]));
    defparam wait_counter_4646_4647_add_4_13.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_13.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_13.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_13.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_11 (.A0(wait_counter[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62748), .COUT(n62749), .S0(n130[9]), 
          .S1(n130[10]));
    defparam wait_counter_4646_4647_add_4_11.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_11.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_11.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_11.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_9 (.A0(wait_counter[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62747), .COUT(n62748), .S0(n130[7]), 
          .S1(n130[8]));
    defparam wait_counter_4646_4647_add_4_9.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_9.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_9.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_9.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_7 (.A0(wait_counter[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62746), .COUT(n62747), .S0(n130[5]), 
          .S1(n130[6]));
    defparam wait_counter_4646_4647_add_4_7.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_7.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_7.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_7.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_5 (.A0(wait_counter[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62745), .COUT(n62746), .S0(n130[3]), 
          .S1(n130[4]));
    defparam wait_counter_4646_4647_add_4_5.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_5.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_5.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_5.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_3 (.A0(wait_counter[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(wait_counter[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n62744), .COUT(n62745), .S0(n130[1]), 
          .S1(n130[2]));
    defparam wait_counter_4646_4647_add_4_3.INIT0 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_3.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_3.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_3.INJECT1_1 = "NO";
    CCU2D wait_counter_4646_4647_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(wait_counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n62744), .S1(n130[0]));
    defparam wait_counter_4646_4647_add_4_1.INIT0 = 16'hF000;
    defparam wait_counter_4646_4647_add_4_1.INIT1 = 16'h0555;
    defparam wait_counter_4646_4647_add_4_1.INJECT1_0 = "NO";
    defparam wait_counter_4646_4647_add_4_1.INJECT1_1 = "NO";
    FD1P3AX div_ce_86_rep_916 (.D(n86), .SP(n142_adj_528), .CK(clock), 
            .Q(n73814));
    defparam div_ce_86_rep_916.GSR = "DISABLED";
    FD1P3AX mul_ce_85_rep_915 (.D(n1442), .SP(n141), .CK(clock), .Q(n73813));
    defparam mul_ce_85_rep_915.GSR = "DISABLED";
    FD1P3AX mul_ce_85_rep_914 (.D(n1442), .SP(n141), .CK(clock), .Q(n73812));
    defparam mul_ce_85_rep_914.GSR = "DISABLED";
    FD1P3AX sub_ce_83_rep_913 (.D(n23885), .SP(n23670), .CK(clock), .Q(n73811));
    defparam sub_ce_83_rep_913.GSR = "DISABLED";
    FD1P3AX sub_ce_83_rep_912 (.D(n23885), .SP(n23670), .CK(clock), .Q(n73810));
    defparam sub_ce_83_rep_912.GSR = "DISABLED";
    LUT4 mux_4234_i1_3_lut (.A(mul_c[0]), .B(div_c[0]), .C(n1148[4]), 
         .Z(n13301[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i1_3_lut.init = 16'hcaca;
    LUT4 i54832_4_lut (.A(n13301[0]), .B(fR1_e3[0]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54832_4_lut.init = 16'h0aca;
    LUT4 i55044_4_lut_rep_911 (.A(wait_counter[17]), .B(n14), .C(n10), 
         .D(wait_counter[21]), .Z(n73809)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i55044_4_lut_rep_911.init = 16'h0001;
    LUT4 mux_4232_i1_3_lut (.A(add_c[0]), .B(sub_c[0]), .C(n1148[2]), 
         .Z(n13267[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i1_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i2_3_lut (.A(mul_c[1]), .B(div_c[1]), .C(n1148[4]), 
         .Z(n13301[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i2_3_lut.init = 16'hcaca;
    LUT4 i54895_4_lut (.A(n13301[1]), .B(fR1_e3[1]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54895_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i2_3_lut (.A(add_c[1]), .B(sub_c[1]), .C(n1148[2]), 
         .Z(n13267[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i2_3_lut.init = 16'hcaca;
    LUT4 mux_4234_i3_3_lut (.A(mul_c[2]), .B(div_c[2]), .C(n1148[4]), 
         .Z(n13301[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i3_3_lut.init = 16'hcaca;
    LUT4 i54893_4_lut (.A(n13301[2]), .B(fR1_e3[2]), .C(n1151), .D(ufl1_e3), 
         .Z(n13369[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i54893_4_lut.init = 16'h0aca;
    LUT4 mux_4232_i3_3_lut (.A(add_c[2]), .B(sub_c[2]), .C(n1148[2]), 
         .Z(n13267[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4232_i3_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n1156), .B(float_alu_mode[0]), .C(\float_alu_mode[1] ), 
         .D(\float_alu_mode[2] ), .Z(n22187)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 mux_4234_i4_3_lut (.A(mul_c[3]), .B(div_c[3]), .C(n1148[4]), 
         .Z(n13301[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4234_i4_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_978 (.A(n1156), .B(float_alu_mode[0]), 
         .C(n1148[4]), .D(\float_alu_mode[2] ), .Z(n86)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_978.init = 16'h0200;
    \fp_add(32,24,8)  fp_sub0 (.clock(clock), .n73811(n73811), .alu_b({alu_b}), 
            .sub_c({sub_c}), .alu_a({alu_a}), .n61(n61), .sub_ce(sub_ce), 
            .\A_int[10] (\A_int[10] ), .\B_int[10] (\B_int[10] ), .n70727(n70727), 
            .\A_int[11] (\A_int[11] ), .\B_int[11] (\B_int[11] ), .\A_int[12] (\A_int[12] ), 
            .\B_int[12] (\B_int[12] ), .n70692(n70692), .\frac[15] (\frac[15] ), 
            .n70693(n70693), .GND_net(GND_net), .diffExpAB({\diffExpAB[8] , 
            Open_58, Open_59, Open_60, Open_61, Open_62, Open_63, 
            Open_64, Open_65}), .n73810(n73810), .n493(n493), .n466(n466), 
            .n70691(n70691), .\efectFracB[13] (\efectFracB[13] ), .\efectFracB[15] (\efectFracB[15] ), 
            .\efectFracB[14] (\efectFracB[14] ));
    \fp_mul(32,24,8)  fp_mul0 (.\B_int[12] (\B_int[12]_adj_2 ), .\B_int[13] (\B_int[13] ), 
            .\B_int[15] (\B_int[15] ), .\B_int[8] (\B_int[8] ), .\A_int[2] (\A_int[2] ), 
            .\A_int[3] (\A_int[3] ), .\A_int[6] (\A_int[6] ), .\A_int[7] (\A_int[7] ), 
            .\A_int[4] (\A_int[4] ), .\A_int[5] (\A_int[5] ), .\B_int[0] (\B_int[0] ), 
            .clock(clock), .n73813(n73813), .alu_b({alu_b}), .\A_int[0] (\A_int[0] ), 
            .alu_a({alu_a}), .\A_int[11] (\A_int[11]_adj_3 ), .\A_int[12] (\A_int[12]_adj_4 ), 
            .\A_int[13] (\A_int[13] ), .\A_int[15] (\A_int[15] ), .\A_int[17] (\A_int[17] ), 
            .\A_int[16] (\A_int[16] ), .\A_int[18] (\A_int[18] ), .\A_int[19] (\A_int[19] ), 
            .\A_int[14] (\A_int[14] ), .n4(n4), .n41520(n41520), .\A_int[1] (\A_int[1] ), 
            .\A_int[10] (\A_int[10]_adj_5 ), .\A_int[9] (\A_int[9] ), .\A_int[22] (\A_int[22] ), 
            .\A_int[21] (\A_int[21] ), .\A_int[8] (\A_int[8] ), .\A_int[20] (\A_int[20] ), 
            .n22310(n22310), .\B_int[11] (\B_int[11]_adj_6 ), .\B_int[14] (\B_int[14] ), 
            .\B_int[10] (\B_int[10]_adj_7 ), .\B_int[9] (\B_int[9] ), .\B_int[19] (\B_int[19] ), 
            .\B_int[18] (\B_int[18] ), .\B_int[20] (\B_int[20] ), .\B_int[21] (\B_int[21] ), 
            .\B_int[7] (\B_int[7] ), .n22437(n22437), .\prod[47] (\prod[47] ), 
            .n66955(n66955), .n67025(n67025), .n67007(n67007), .n41808(n41808), 
            .\prod[45] (\prod[45] ), .\prod[46] (\prod[46] ), .\prod[28] (\prod[28] ), 
            .\prod[33] (\prod[33] ), .\prod[40] (\prod[40] ), .\prod[22] (\prod[22] ), 
            .\prod[24] (\prod[24] ), .\prod[25] (\prod[25] ), .\prod[23] (\prod[23] ), 
            .\prod[26] (\prod[26] ), .\prod[41] (\prod[41] ), .\prod[34] (\prod[34] ), 
            .\prod[37] (\prod[37] ), .\prod[27] (\prod[27] ), .\prod[39] (\prod[39] ), 
            .\prod[29] (\prod[29] ), .\prod[35] (\prod[35] ), .\prod[36] (\prod[36] ), 
            .\prod[31] (\prod[31] ), .\prod[32] (\prod[32] ), .\prod[43] (\prod[43] ), 
            .\prod[30] (\prod[30] ), .\prod[38] (\prod[38] ), .\prod[42] (\prod[42] ), 
            .\prod[44] (\prod[44] ), .n42939(n42939), .n42941(n42941), 
            .n25571(n25571), .n73812(n73812), .n42934(n42934), .mul_c({mul_c}), 
            .GND_net(GND_net), .\frac_norm[20] (\frac_norm[20] ), .\frac_norm[16] (\frac_norm[16] ), 
            .\frac_norm[14] (\frac_norm[14] ), .\frac_norm[15] (\frac_norm[15] ), 
            .\frac_norm[12] (\frac_norm[12] ), .\frac_norm[13] (\frac_norm[13] ), 
            .\frac_norm[10] (\frac_norm[10] ), .\frac_norm[11] (\frac_norm[11] ), 
            .\frac_norm[8] (\frac_norm[8] ), .n15(n15), .\B_int[17] (\B_int[17] ), 
            .\B_int[16] (\B_int[16] ), .\B_int[22] (\B_int[22] ), .\frac_norm[7] (\frac_norm[7] ), 
            .n25583(n25583), .n984({n984}), .\B_int[3] (\B_int[3] ), .\B_int[1] (\B_int[1] ), 
            .\B_int[2] (\B_int[2] ), .\frac_norm[4] (\frac_norm[4] ), .\frac_norm[5] (\frac_norm[5] ), 
            .\frac_norm[3] (\frac_norm[3] ), .\frac_norm[2] (\frac_norm[2] ), 
            .exp_final({exp_final}), .\FP_Z_int[22] (\FP_Z_int[22] ), .mul_ce(mul_ce), 
            .\B_int[6] (\B_int[6] ), .\B_int[5] (\B_int[5] ), .\B_int[4] (\B_int[4] ), 
            .n6(n6), .\prod[21] (\prod[21] ));
    \fp_exp_clk(8,23)  fp_exp_clk0 (.clock(clock), .fR1_e3({Open_66, Open_67, 
            Open_68, Open_69, Open_70, Open_71, Open_72, Open_73, 
            Open_74, Open_75, Open_76, Open_77, Open_78, Open_79, 
            Open_80, Open_81, Open_82, Open_83, Open_84, Open_85, 
            Open_86, Open_87, Open_88, fR1_e3[0]}), .GND_net(GND_net), 
            .ufl1_e3(ufl1_e3), .\fR1_e3[22] (fR1_e3[22]), .\fR1_e3[21] (fR1_e3[21]), 
            .\fR1_e3[20] (fR1_e3[20]), .\fR1_e3[19] (fR1_e3[19]), .\fR1_e3[18] (fR1_e3[18]), 
            .\fR1_e3[17] (fR1_e3[17]), .\fR1_e3[16] (fR1_e3[16]), .\fR1_e3[15] (fR1_e3[15]), 
            .\fR1_e3[14] (fR1_e3[14]), .\fR1_e3[13] (fR1_e3[13]), .\fR1_e3[12] (fR1_e3[12]), 
            .\fR1_e3[11] (fR1_e3[11]), .\fR1_e3[10] (fR1_e3[10]), .\fR1_e3[9] (fR1_e3[9]), 
            .\fR1_e3[8] (fR1_e3[8]), .\fR1_e3[7] (fR1_e3[7]), .\fR1_e3[6] (fR1_e3[6]), 
            .\fR1_e3[5] (fR1_e3[5]), .\fR1_e3[4] (fR1_e3[4]), .\fR1_e3[3] (fR1_e3[3]), 
            .\fR1_e3[2] (fR1_e3[2]), .\fR1_e3[1] (fR1_e3[1]), .\eR_e3[7] (eR_e3[7]), 
            .\eR_e3[5] (eR_e3[5]), .\eR_e3[6] (eR_e3[6]), .\eR_e3[3] (eR_e3[3]), 
            .\eR_e3[4] (eR_e3[4]), .\eR_e3[1] (eR_e3[1]), .\eR_e3[2] (eR_e3[2]), 
            .\eR_e3[0] (eR_e3[0]), .\mXs_0[24] (mXs_0[24]), .\exp_a[0] (exp_a[0]), 
            .\exp_a[1] (exp_a[1]), .\exp_a[2] (exp_a[2]), .\exp_a[3] (exp_a[3]), 
            .\exp_a[4] (exp_a[4]), .\exp_a[5] (exp_a[5]), .\exp_a[6] (exp_a[6]), 
            .\exp_a[7] (exp_a[7]), .\exp_a[8] (exp_a[8]), .\exp_a[9] (exp_a[9]), 
            .\exp_a[10] (exp_a[10]), .\exp_a[11] (exp_a[11]), .\exp_a[12] (exp_a[12]), 
            .\exp_a[13] (exp_a[13]), .\exp_a[14] (exp_a[14]), .\exp_a[15] (exp_a[15]), 
            .\exp_a[16] (exp_a[16]), .\exp_a[17] (exp_a[17]), .\exp_a[18] (exp_a[18]), 
            .\exp_a[19] (exp_a[19]), .\exp_a[20] (exp_a[20]), .\exp_a[21] (exp_a[21]), 
            .\exp_a[22] (exp_a[22]), .\exp_a[30] (exp_a[30]), .\exp_a[28] (exp_a[28]), 
            .\exp_a[29] (exp_a[29]), .\exp_a[26] (exp_a[26]), .\exp_a[27] (exp_a[27]), 
            .\exp_a[24] (exp_a[24]), .\exp_a[25] (exp_a[25]), .\exp_a[23] (exp_a[23]), 
            .VCC_net(VCC_net), .\buf_x[89] (\buf_x[89] ), .\buf_x[87] (\buf_x[87] ), 
            .\buf_x[88] (\buf_x[88] ), .\buf_x[85] (\buf_x[85] ), .\buf_x[86] (\buf_x[86] ), 
            .\buf_x[83] (\buf_x[83] ), .\buf_x[84] (\buf_x[84] ), .\buf_r[89] (\buf_r[89] ), 
            .\buf_r[87] (\buf_r[87] ), .\buf_r[88] (\buf_r[88] ), .\buf_r[85] (\buf_r[85] ), 
            .\buf_r[86] (\buf_r[86] ), .\buf_r[83] (\buf_r[83] ), .\buf_r[84] (\buf_r[84] ), 
            .\exp_a[32] (exp_a[32]));
    \fp_div(32,24,8)  fp_div0 (.GND_net(GND_net), .clock(clock), .n73815(n73815), 
            .alu_b({alu_b}), .alu_a({alu_a}), .div_c({div_c}), .div_ce(div_ce), 
            .n73814(n73814));
    \fp_add(32,24,8)_U28  fp_add0 (.add_c({add_c}), .clock(clock), .n73804(n73804), 
            .\A_int[11] (\A_int[11]_adj_8 ), .\B_int[11] (\B_int[11]_adj_9 ), 
            .\A_int[10] (\A_int[10]_adj_10 ), .\B_int[10] (\B_int[10]_adj_11 ), 
            .\A_int[13] (\A_int[13]_adj_12 ), .\B_int[13] (\B_int[13]_adj_13 ), 
            .\A_int[12] (\A_int[12]_adj_14 ), .\B_int[12] (\B_int[12]_adj_15 ), 
            .add_ce(add_ce), .\A_int[17] (\A_int[17]_adj_16 ), .\B_int[17] (\B_int[17]_adj_17 ), 
            .alu_b({alu_b}), .\A_int[16] (\A_int[16]_adj_18 ), .\B_int[16] (\B_int[16]_adj_19 ), 
            .alu_a({alu_a}), .\A_int[18] (\A_int[18]_adj_20 ), .\B_int[18] (\B_int[18]_adj_21 ), 
            .GND_net(GND_net), .\A_int[2] (\A_int[2]_adj_22 ), .\B_int[2] (\B_int[2]_adj_23 ), 
            .\B_int[3] (\B_int[3]_adj_24 ), .\A_int[9] (\A_int[9]_adj_25 ), 
            .\A_int[7] (\A_int[7]_adj_26 ), .\A_int[4] (\A_int[4]_adj_27 ), 
            .\A_int[3] (\A_int[3]_adj_28 ), .\B_int[9] (\B_int[9]_adj_29 ), 
            .\B_int[7] (\B_int[7]_adj_30 ), .\B_int[4] (\B_int[4]_adj_31 ), 
            .diffExpAB({\diffExpAB[8]_adj_32 , Open_89, Open_90, Open_91, 
            Open_92, Open_93, Open_94, Open_95, Open_96}), .add_enable(add_enable), 
            .\diffExp[4] (\diffExp[4] ), .n73803(n73803), .n70835(n70835), 
            .n70834(n70834), .n70833(n70833), .\efectFracB[21] (\efectFracB[21] ), 
            .\efectFracB[20] (\efectFracB[20] ), .\efectFracB[19] (\efectFracB[19] ), 
            .\efectFracB[15] (\efectFracB[15]_adj_33 ), .\efectFracB[16] (\efectFracB[16] ), 
            .n19214(n19214), .n28(n28), .n70771(n70771), .n9(n9), .\efectFracB[14] (\efectFracB[14]_adj_34 ), 
            .\efectFracB[7] (\efectFracB[7] ), .\efectFracB[5] (\efectFracB[5] ), 
            .\efectFracB[12] (\efectFracB[12] ), .n70820(n70820), .\efectFracB[13] (\efectFracB[13]_adj_35 ), 
            .n27(n27), .n70740(n70740), .n55(n55));
    
endmodule
//
// Verilog Description of module \fp_add(32,24,8) 
//

module \fp_add(32,24,8)  (clock, n73811, alu_b, sub_c, alu_a, n61, 
            sub_ce, \A_int[10] , \B_int[10] , n70727, \A_int[11] , 
            \B_int[11] , \A_int[12] , \B_int[12] , n70692, \frac[15] , 
            n70693, GND_net, diffExpAB, n73810, n493, n466, n70691, 
            \efectFracB[13] , \efectFracB[15] , \efectFracB[14] );
    input clock;
    input n73811;
    input [31:0]alu_b;
    output [31:0]sub_c;
    input [31:0]alu_a;
    output n61;
    input sub_ce;
    output \A_int[10] ;
    output \B_int[10] ;
    output n70727;
    output \A_int[11] ;
    output \B_int[11] ;
    output \A_int[12] ;
    output \B_int[12] ;
    input n70692;
    input \frac[15] ;
    output n70693;
    input GND_net;
    output [8:0]diffExpAB;
    input n73810;
    output n493;
    output n466;
    input n70691;
    input \efectFracB[13] ;
    input \efectFracB[15] ;
    input \efectFracB[14] ;
    
    wire [31:0]A_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(54[11:16])
    wire [31:0]B_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(55[11:16])
    wire [4:0]leadZerosBin;   // c:/users/yisong/documents/new/mlp/fp_leading_zeros_and_shift.vhd(25[11:23])
    wire [27:0]subBAExpEq;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(73[11:21])
    wire isSUB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(71[11:16])
    wire [27:0]fracAlign_int;   // c:/users/yisong/documents/new/mlp/right_shifter.vhd(21[11:24])
    wire [31:0]FP_Z_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(106[11:19])
    wire [27:0]frac_Norm1;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(97[17:27])
    wire [27:0]addSubAB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(69[18:26])
    wire [22:0]frac_Norm2;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(98[11:21])
    wire [27:0]frac;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(97[11:15])
    wire [8:0]efectExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(65[11:19])
    wire [27:0]frac_add_Norm1;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(70[11:25])
    wire [27:0]frac_sub_Norm1;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(74[11:25])
    wire sign;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(75[11:15])
    wire [8:0]diffExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[33:40])
    wire [8:0]diffExpAB_c;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[11:20])
    wire [27:0]efectFracB_align;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(67[35:51])
    wire expA_FF;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(56[11:18])
    wire expB_FF;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(56[20:27])
    wire [8:0]diffExpBA;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[22:31])
    
    wire n41452, n73796, n41448, n41450, n448, n70738, n7, n21707, 
        n21703, n21701, n15583, n21731, n21673, n21697, n15599, 
        n21741, n21721, n21723, n21729, n21743, n21733, n21735, 
        n21727, n70133, n70134, n41445, n41499, n21739, n21737, 
        n40001, n62960, n53, n70612, n70837, n70634, n70721, n66873, 
        n43011, n41366, n41374, n41382, n24092;
    wire [22:0]n10672;
    
    wire n41384, n41386, n41388, n41390, n41392, n41394, n41396;
    wire [27:0]n451;
    wire [27:0]n480;
    
    wire n41404, n41406, n41418, n41420, n41441, n41443, n41501, 
        n39997, n39999, n70729, n770, n769, n768, n767, n766, 
        n765, n764, n763;
    wire [7:0]n8351;
    
    wire n103, n73797, n70635, n70639;
    wire [27:0]n243;
    
    wire n66231, n731, n41446, n70067, n70618, n4, n70620, n70782, 
        n70677, n70680, n70681, n17520, n66711, n70617, n18;
    wire [27:0]n330;
    
    wire n66709, n79, n70683;
    wire [27:0]n301;
    
    wire n9, n11, n70688, n70687, n70689, n41774, n7_adj_497, 
        n73798, n70132, n70131, n60994, n60993, n61566, n61565, 
        n70717, n73142, n73141, n67674, n73140, n41776, n21699, 
        n61564, n73139, n70676, n70709, n70763, n41584, n21717, 
        n70718, n15, n70734, n21719, n66912, n21725, n66898, n21715, 
        n66185, n9_adj_498, n14, n10, n61563, n61562, n61561, 
        n61560, n61559, n61558, n61557, n61556, n70626, n66825, 
        n70625, n70698, n73799, n70710, n41732, n61839, n61838, 
        n66221, n61555, n70699, n70704, n61837, n61836, n61835, 
        n61834, n61833, n61832, n61831, n61830, n61829, n61553, 
        n61828, n61827, n61826, n61552, n61551, n61550, n10_adj_499, 
        n14_adj_500, n10_adj_501, n14_adj_502, n44, n34, n48, n41, 
        n40, n31, n32, n50, n45, n39, n93, n10_adj_503, n16, 
        n15_adj_504, n22573, n66199, n4_adj_505, n61548, n61547, 
        n61546, n61545, n22515, n70658, n70647, n61544, n61543, 
        n41812, n70690, n28, n38, n24, n36, n42, n61542, n32_adj_506, 
        n40_adj_507, n44_adj_508, n31_adj_509, n10_adj_510, n14_adj_511, 
        n9_adj_512, n61541, n41444, n41498, n40000, n61540, n28_adj_513, 
        n38_adj_514, n24_adj_515, n36_adj_516, n42_adj_517, n41365, 
        n41373, n41381, n32_adj_518, n40_adj_519, n41383, n44_adj_520, 
        n31_adj_521, n41385, n61539, n41391, n61538, n63641, n41393, 
        n41395, n41403, n41405, n41417, n41500, n41442, n41389, 
        n41440, n39998, n39996, n41419, n41387, n39_adj_522, n41_adj_523, 
        n30, n45_adj_524, n37, n44_adj_525, n33, n34_adj_526, n48_adj_527, 
        n43, n574, n62172, n62171, n62170, n62169, n61621, n61620, 
        n61619, n61618;
    wire [27:0]n272;
    
    wire n66493;
    
    LUT4 i29857_2_lut_3_lut (.A(A_int[31]), .B(B_int[31]), .C(leadZerosBin[1]), 
         .Z(n41452)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam i29857_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i29853_2_lut_3_lut (.A(A_int[31]), .B(B_int[31]), .C(n73796), 
         .Z(n41448)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam i29853_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i29855_2_lut_3_lut (.A(A_int[31]), .B(B_int[31]), .C(leadZerosBin[2]), 
         .Z(n41450)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam i29855_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i2_3_lut_rep_768_4_lut (.A(A_int[31]), .B(B_int[31]), .C(subBAExpEq[27]), 
         .D(n448), .Z(n70738)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B+(C+!(D)))) */ ;
    defparam i2_3_lut_rep_768_4_lut.init = 16'hf6ff;
    LUT4 i10009_1_lut_2_lut (.A(A_int[31]), .B(B_int[31]), .Z(isSUB)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i10009_1_lut_2_lut.init = 16'h9999;
    LUT4 i1_3_lut_4_lut (.A(A_int[31]), .B(B_int[31]), .C(n7), .D(fracAlign_int[4]), 
         .Z(n21707)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_900 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[3]), .Z(n21703)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_900.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_901 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[6]), .Z(n21701)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_901.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_902 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[5]), .Z(n15583)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_902.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_903 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[8]), .Z(n21731)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_903.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_904 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[7]), .Z(n21673)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_904.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_905 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[10]), .Z(n21697)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_905.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_906 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[9]), .Z(n15599)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_906.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_907 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[12]), .Z(n21741)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_907.init = 16'h6966;
    FD1P3AX B_int_i0_i0 (.D(alu_b[0]), .SP(n73811), .CK(clock), .Q(B_int[0]));
    defparam B_int_i0_i0.GSR = "DISABLED";
    FD1P3AX FP_Z_i0_i0 (.D(FP_Z_int[0]), .SP(n73811), .CK(clock), .Q(sub_c[0]));
    defparam FP_Z_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_908 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[14]), .Z(n21721)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_908.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_909 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[13]), .Z(n21723)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_909.init = 16'h6966;
    FD1P3AX A_int_i0_i0 (.D(alu_a[0]), .SP(n73811), .CK(clock), .Q(A_int[0]));
    defparam A_int_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_910 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[16]), .Z(n21729)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_910.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_911 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[15]), .Z(n21743)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_911.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_912 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[18]), .Z(n21733)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_912.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_913 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[17]), .Z(n21735)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_913.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_914 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[20]), .Z(n21727)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_914.init = 16'h6966;
    LUT4 n70134_bdd_3_lut_4_lut (.A(A_int[31]), .B(B_int[31]), .C(n70133), 
         .D(n70134), .Z(frac_Norm1[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n70134_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 i29850_3_lut (.A(A_int[17]), .B(B_int[17]), .C(n61), .Z(n41445)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29850_3_lut.init = 16'hacac;
    LUT4 i29904_3_lut (.A(A_int[18]), .B(B_int[18]), .C(n61), .Z(n41499)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29904_3_lut.init = 16'hacac;
    LUT4 i1_3_lut_4_lut_adj_915 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[21]), .Z(n21739)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_915.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_916 (.A(A_int[31]), .B(B_int[31]), .C(n7), 
         .D(fracAlign_int[22]), .Z(n21737)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_916.init = 16'h6966;
    LUT4 i28408_3_lut (.A(A_int[22]), .B(B_int[22]), .C(n61), .Z(n40001)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i28408_3_lut.init = 16'hacac;
    LUT4 i28149_3_lut_rep_642_4_lut (.A(A_int[31]), .B(B_int[31]), .C(n62960), 
         .D(n53), .Z(n70612)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B+(C (D)))) */ ;
    defparam i28149_3_lut_rep_642_4_lut.init = 16'hf666;
    LUT4 i1_2_lut_rep_867 (.A(A_int[31]), .B(B_int[31]), .Z(n70837)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_867.init = 16'h6666;
    LUT4 i2_3_lut_4_lut (.A(n70634), .B(n70721), .C(addSubAB[2]), .D(n66873), 
         .Z(n43011)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 i29773_3_lut (.A(A_int[1]), .B(B_int[1]), .C(n61), .Z(n41366)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29773_3_lut.init = 16'hacac;
    LUT4 i29781_3_lut (.A(A_int[2]), .B(B_int[2]), .C(n61), .Z(n41374)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29781_3_lut.init = 16'hacac;
    LUT4 i29789_3_lut (.A(A_int[3]), .B(B_int[3]), .C(n61), .Z(n41382)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29789_3_lut.init = 16'hacac;
    FD1P3IX FP_Z_i0_i1 (.D(n10672[1]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[1]));
    defparam FP_Z_i0_i1.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i2 (.D(n10672[2]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[2]));
    defparam FP_Z_i0_i2.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i3 (.D(n10672[3]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[3]));
    defparam FP_Z_i0_i3.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i4 (.D(n10672[4]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[4]));
    defparam FP_Z_i0_i4.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i5 (.D(n10672[5]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[5]));
    defparam FP_Z_i0_i5.GSR = "DISABLED";
    LUT4 i29791_3_lut (.A(A_int[4]), .B(B_int[4]), .C(n61), .Z(n41384)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29791_3_lut.init = 16'hacac;
    LUT4 i29793_3_lut (.A(A_int[5]), .B(B_int[5]), .C(n61), .Z(n41386)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29793_3_lut.init = 16'hacac;
    FD1P3IX FP_Z_i0_i6 (.D(n10672[6]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[6]));
    defparam FP_Z_i0_i6.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i7 (.D(n10672[7]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[7]));
    defparam FP_Z_i0_i7.GSR = "DISABLED";
    LUT4 i29795_3_lut (.A(A_int[6]), .B(B_int[6]), .C(n61), .Z(n41388)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29795_3_lut.init = 16'hacac;
    LUT4 i29797_3_lut (.A(A_int[7]), .B(B_int[7]), .C(n61), .Z(n41390)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29797_3_lut.init = 16'hacac;
    LUT4 i29799_3_lut (.A(A_int[8]), .B(B_int[8]), .C(n61), .Z(n41392)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29799_3_lut.init = 16'hacac;
    LUT4 i29801_3_lut (.A(A_int[9]), .B(B_int[9]), .C(n61), .Z(n41394)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29801_3_lut.init = 16'hacac;
    LUT4 i29803_3_lut (.A(\A_int[10] ), .B(\B_int[10] ), .C(n61), .Z(n41396)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29803_3_lut.init = 16'hacac;
    LUT4 mux_52_i4_3_lut (.A(A_int[0]), .B(n451[3]), .C(n70727), .Z(n480[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i4_3_lut.init = 16'hcaca;
    LUT4 i29811_3_lut (.A(\A_int[11] ), .B(\B_int[11] ), .C(n61), .Z(n41404)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29811_3_lut.init = 16'hacac;
    LUT4 i29813_3_lut (.A(\A_int[12] ), .B(\B_int[12] ), .C(n61), .Z(n41406)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29813_3_lut.init = 16'hacac;
    LUT4 i29825_3_lut (.A(A_int[13]), .B(B_int[13]), .C(n61), .Z(n41418)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29825_3_lut.init = 16'hacac;
    LUT4 i29827_3_lut (.A(A_int[14]), .B(B_int[14]), .C(n61), .Z(n41420)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29827_3_lut.init = 16'hacac;
    LUT4 i29846_3_lut (.A(A_int[15]), .B(B_int[15]), .C(n61), .Z(n41441)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29846_3_lut.init = 16'hacac;
    LUT4 i29848_3_lut (.A(A_int[16]), .B(B_int[16]), .C(n61), .Z(n41443)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29848_3_lut.init = 16'hacac;
    LUT4 i29906_3_lut (.A(A_int[19]), .B(B_int[19]), .C(n61), .Z(n41501)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29906_3_lut.init = 16'hacac;
    LUT4 i28404_3_lut (.A(A_int[20]), .B(B_int[20]), .C(n61), .Z(n39997)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i28404_3_lut.init = 16'hacac;
    LUT4 i28406_3_lut (.A(A_int[21]), .B(B_int[21]), .C(n61), .Z(n39999)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i28406_3_lut.init = 16'hacac;
    FD1P3IX FP_Z_i0_i8 (.D(n10672[8]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[8]));
    defparam FP_Z_i0_i8.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i9 (.D(n10672[9]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[9]));
    defparam FP_Z_i0_i9.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i10 (.D(n10672[10]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[10]));
    defparam FP_Z_i0_i10.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i11 (.D(n10672[11]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[11]));
    defparam FP_Z_i0_i11.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i12 (.D(n10672[12]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[12]));
    defparam FP_Z_i0_i12.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i13 (.D(n10672[13]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[13]));
    defparam FP_Z_i0_i13.GSR = "DISABLED";
    LUT4 mux_3772_i1_4_lut (.A(frac_Norm2[0]), .B(frac[3]), .C(n70729), 
         .D(n70612), .Z(n10672[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i1_4_lut.init = 16'hcac0;
    FD1P3IX FP_Z_i0_i14 (.D(n10672[14]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[14]));
    defparam FP_Z_i0_i14.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i15 (.D(n10672[15]), .SP(sub_ce), .CD(n24092), .CK(clock), 
            .Q(sub_c[15]));
    defparam FP_Z_i0_i15.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i16 (.D(n10672[16]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[16]));
    defparam FP_Z_i0_i16.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i17 (.D(n10672[17]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[17]));
    defparam FP_Z_i0_i17.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i18 (.D(n10672[18]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[18]));
    defparam FP_Z_i0_i18.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i19 (.D(n10672[19]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[19]));
    defparam FP_Z_i0_i19.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i20 (.D(n10672[20]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[20]));
    defparam FP_Z_i0_i20.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i21 (.D(n10672[21]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[21]));
    defparam FP_Z_i0_i21.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i22 (.D(n10672[22]), .SP(n73811), .CD(n24092), .CK(clock), 
            .Q(sub_c[22]));
    defparam FP_Z_i0_i22.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i23 (.D(n770), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[23]));
    defparam FP_Z_i0_i23.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i24 (.D(n769), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[24]));
    defparam FP_Z_i0_i24.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i25 (.D(n768), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[25]));
    defparam FP_Z_i0_i25.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i26 (.D(n767), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[26]));
    defparam FP_Z_i0_i26.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i27 (.D(n766), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[27]));
    defparam FP_Z_i0_i27.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i28 (.D(n765), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[28]));
    defparam FP_Z_i0_i28.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i29 (.D(n764), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[29]));
    defparam FP_Z_i0_i29.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i30 (.D(n763), .SP(n73811), .PD(n24092), .CK(clock), 
            .Q(sub_c[30]));
    defparam FP_Z_i0_i30.GSR = "DISABLED";
    LUT4 i110_4_lut (.A(n8351[7]), .B(efectExp[7]), .C(n70729), .D(n103), 
         .Z(n763)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i110_4_lut.init = 16'hcac0;
    LUT4 i28184_2_lut_4_lut (.A(n73797), .B(n70635), .C(n70639), .D(frac[12]), 
         .Z(n243[12])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28184_2_lut_4_lut.init = 16'h8000;
    LUT4 i28186_2_lut_4_lut (.A(n73797), .B(n70635), .C(n70639), .D(frac[10]), 
         .Z(n243[10])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28186_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut (.A(n10672[0]), .B(n66231), .C(n731), .Z(FP_Z_int[0])) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i1_3_lut.init = 16'hcece;
    LUT4 i29851_2_lut_4_lut (.A(n73797), .B(n70635), .C(n70639), .D(n70837), 
         .Z(n41446)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i29851_2_lut_4_lut.init = 16'hff7f;
    LUT4 n1_bdd_2_lut_55850_rep_648_4_lut (.A(n73797), .B(n70635), .C(n70639), 
         .D(n70067), .Z(n70618)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam n1_bdd_2_lut_55850_rep_648_4_lut.init = 16'h8000;
    LUT4 i111_4_lut (.A(n8351[6]), .B(efectExp[6]), .C(n70729), .D(n103), 
         .Z(n764)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i111_4_lut.init = 16'hcac0;
    LUT4 i15319_4_lut (.A(n8351[5]), .B(efectExp[5]), .C(n70729), .D(n103), 
         .Z(n765)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i15319_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_4_lut (.A(n73797), .B(n70635), .C(n70639), .D(frac[3]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i28183_2_lut_4_lut (.A(n73797), .B(n70635), .C(n70639), .D(n70692), 
         .Z(n243[13])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28183_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_650_4_lut (.A(n73797), .B(n70635), .C(n70639), .D(efectExp[4]), 
         .Z(n70620)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i1_2_lut_rep_650_4_lut.init = 16'h7f80;
    LUT4 i15324_4_lut (.A(n8351[4]), .B(efectExp[4]), .C(n70729), .D(n103), 
         .Z(n766)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i15324_4_lut.init = 16'hcac0;
    LUT4 i114_4_lut (.A(n8351[3]), .B(n70782), .C(n70729), .D(n103), 
         .Z(n767)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i114_4_lut.init = 16'hcac0;
    LUT4 i115_4_lut (.A(n8351[2]), .B(efectExp[2]), .C(n70729), .D(n103), 
         .Z(n768)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i115_4_lut.init = 16'hcac0;
    LUT4 i116_4_lut (.A(n8351[1]), .B(efectExp[1]), .C(n70729), .D(n103), 
         .Z(n769)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i116_4_lut.init = 16'hcac0;
    LUT4 i117_4_lut (.A(n8351[0]), .B(efectExp[0]), .C(n70729), .D(n103), 
         .Z(n770)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i117_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i23_4_lut (.A(frac_Norm2[22]), .B(n70677), .C(n70729), 
         .D(n70612), .Z(n10672[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i23_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i22_4_lut (.A(frac_Norm2[21]), .B(n70680), .C(n70729), 
         .D(n70612), .Z(n10672[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i22_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i21_4_lut (.A(frac_Norm2[20]), .B(n70681), .C(n70729), 
         .D(n70612), .Z(n10672[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i21_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut (.A(frac_Norm1[3]), .B(addSubAB[0]), .C(n17520), .D(leadZerosBin[1]), 
         .Z(n66711)) /* synthesis lut_function=(A+!((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'haaae;
    LUT4 i1_4_lut_adj_917 (.A(addSubAB[1]), .B(n70617), .C(leadZerosBin[2]), 
         .D(leadZerosBin[1]), .Z(n18)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_917.init = 16'h0002;
    LUT4 i31626_4_lut (.A(n43011), .B(addSubAB[0]), .C(leadZerosBin[1]), 
         .D(n17520), .Z(n330[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i31626_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_918 (.A(frac_add_Norm1[2]), .B(frac_Norm1[3]), .C(n70721), 
         .D(n66709), .Z(n79)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_918.init = 16'ha888;
    LUT4 mux_3772_i20_4_lut (.A(frac_Norm2[19]), .B(n70683), .C(n70729), 
         .D(n70612), .Z(n10672[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i20_4_lut.init = 16'hcac0;
    LUT4 i31628_3_lut (.A(n301[4]), .B(n43011), .C(leadZerosBin[1]), .Z(n330[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31628_3_lut.init = 16'hcaca;
    LUT4 i31633_3_lut (.A(n301[6]), .B(n301[4]), .C(leadZerosBin[1]), 
         .Z(n330[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31633_3_lut.init = 16'hcaca;
    LUT4 i9_3_lut (.A(n301[8]), .B(n301[6]), .C(leadZerosBin[1]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9_3_lut.init = 16'hcaca;
    LUT4 i16_3_lut (.A(n330[9]), .B(n9), .C(leadZerosBin[0]), .Z(frac_sub_Norm1[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i16_3_lut.init = 16'hcaca;
    LUT4 i10_3_lut (.A(n9), .B(n330[7]), .C(leadZerosBin[0]), .Z(frac_sub_Norm1[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i10_3_lut.init = 16'hcaca;
    LUT4 mux_3772_i19_4_lut (.A(frac_Norm2[18]), .B(frac[21]), .C(n70729), 
         .D(n70612), .Z(n10672[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i19_4_lut.init = 16'hcac0;
    LUT4 i11_3_lut (.A(n301[10]), .B(n301[8]), .C(leadZerosBin[1]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 mux_3772_i18_4_lut (.A(frac_Norm2[17]), .B(n70688), .C(n70729), 
         .D(n70612), .Z(n10672[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i18_4_lut.init = 16'hcac0;
    LUT4 i14_3_lut (.A(n330[11]), .B(n11), .C(leadZerosBin[0]), .Z(frac_sub_Norm1[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14_3_lut.init = 16'hcaca;
    LUT4 mux_3772_i17_4_lut (.A(frac_Norm2[16]), .B(n70687), .C(n70729), 
         .D(n70612), .Z(n10672[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i17_4_lut.init = 16'hcac0;
    LUT4 i12_3_lut (.A(n11), .B(n330[9]), .C(leadZerosBin[0]), .Z(frac_sub_Norm1[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12_3_lut.init = 16'hcaca;
    LUT4 mux_3772_i16_4_lut (.A(frac_Norm2[15]), .B(frac[18]), .C(n70729), 
         .D(n70612), .Z(n10672[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i16_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i15_4_lut (.A(frac_Norm2[14]), .B(n70689), .C(n70729), 
         .D(n70612), .Z(n10672[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i15_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i14_4_lut (.A(frac_Norm2[13]), .B(frac[16]), .C(n70729), 
         .D(n70612), .Z(n10672[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i14_4_lut.init = 16'hcac0;
    LUT4 i7_4_lut (.A(n70634), .B(n301[10]), .C(leadZerosBin[1]), .D(n41774), 
         .Z(n7_adj_497)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i7_4_lut.init = 16'hcac0;
    LUT4 i8_3_lut (.A(n330[13]), .B(n7_adj_497), .C(leadZerosBin[0]), 
         .Z(frac_sub_Norm1[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i8_3_lut.init = 16'hcaca;
    LUT4 i6_3_lut (.A(n7_adj_497), .B(n330[11]), .C(leadZerosBin[0]), 
         .Z(frac_sub_Norm1[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i6_3_lut.init = 16'hcaca;
    LUT4 mux_3772_i13_4_lut (.A(frac_Norm2[12]), .B(\frac[15] ), .C(n70729), 
         .D(n70612), .Z(n10672[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i13_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i12_4_lut (.A(frac_Norm2[11]), .B(n70693), .C(n70729), 
         .D(n70612), .Z(n10672[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i12_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i11_4_lut (.A(frac_Norm2[10]), .B(n70692), .C(n70729), 
         .D(n70612), .Z(n10672[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i11_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i10_4_lut (.A(frac_Norm2[9]), .B(frac[12]), .C(n70729), 
         .D(n70612), .Z(n10672[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i10_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i9_4_lut (.A(frac_Norm2[8]), .B(n73798), .C(n70729), 
         .D(n70612), .Z(n10672[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i9_4_lut.init = 16'hcac0;
    PFUMX i55875 (.BLUT(n70132), .ALUT(n70131), .C0(n70729), .Z(n70133));
    LUT4 n6_bdd_3_lut_55874 (.A(B_int[0]), .B(n61), .C(A_int[0]), .Z(n70131)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6_bdd_3_lut_55874.init = 16'he2e2;
    CCU2D equal_48_8 (.A0(B_int[24]), .B0(A_int[24]), .C0(B_int[23]), 
          .D0(A_int[23]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n60994), .S1(n448));
    defparam equal_48_8.INIT0 = 16'h9009;
    defparam equal_48_8.INIT1 = 16'hFFFF;
    defparam equal_48_8.INJECT1_0 = "YES";
    defparam equal_48_8.INJECT1_1 = "NO";
    CCU2D equal_48_7 (.A0(B_int[28]), .B0(A_int[28]), .C0(B_int[27]), 
          .D0(A_int[27]), .A1(B_int[26]), .B1(A_int[26]), .C1(B_int[25]), 
          .D1(A_int[25]), .CIN(n60993), .COUT(n60994));
    defparam equal_48_7.INIT0 = 16'h9009;
    defparam equal_48_7.INIT1 = 16'h9009;
    defparam equal_48_7.INJECT1_0 = "YES";
    defparam equal_48_7.INJECT1_1 = "YES";
    CCU2D equal_48_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(B_int[30]), .B1(A_int[30]), .C1(B_int[29]), .D1(A_int[29]), 
          .COUT(n60993));
    defparam equal_48_0.INIT0 = 16'hF000;
    defparam equal_48_0.INIT1 = 16'h9009;
    defparam equal_48_0.INJECT1_0 = "NO";
    defparam equal_48_0.INJECT1_1 = "YES";
    CCU2D sub_214_add_2_25 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61566), .S0(subBAExpEq[26]), .S1(subBAExpEq[27]));
    defparam sub_214_add_2_25.INIT0 = 16'h0fff;
    defparam sub_214_add_2_25.INIT1 = 16'hffff;
    defparam sub_214_add_2_25.INJECT1_0 = "NO";
    defparam sub_214_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_23 (.A0(B_int[21]), .B0(A_int[21]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[22]), .B1(A_int[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61565), .COUT(n61566), .S0(subBAExpEq[24]), 
          .S1(subBAExpEq[25]));
    defparam sub_214_add_2_23.INIT0 = 16'h5999;
    defparam sub_214_add_2_23.INIT1 = 16'h5999;
    defparam sub_214_add_2_23.INJECT1_0 = "NO";
    defparam sub_214_add_2_23.INJECT1_1 = "NO";
    FD1P3AX A_int_i0_i31 (.D(alu_a[31]), .SP(n73811), .CK(clock), .Q(A_int[31]));
    defparam A_int_i0_i31.GSR = "DISABLED";
    FD1P3AX A_int_i0_i30 (.D(alu_a[30]), .SP(n73811), .CK(clock), .Q(A_int[30]));
    defparam A_int_i0_i30.GSR = "DISABLED";
    FD1P3AX A_int_i0_i29 (.D(alu_a[29]), .SP(n73811), .CK(clock), .Q(A_int[29]));
    defparam A_int_i0_i29.GSR = "DISABLED";
    FD1P3AX A_int_i0_i28 (.D(alu_a[28]), .SP(n73811), .CK(clock), .Q(A_int[28]));
    defparam A_int_i0_i28.GSR = "DISABLED";
    FD1P3AX A_int_i0_i27 (.D(alu_a[27]), .SP(n73811), .CK(clock), .Q(A_int[27]));
    defparam A_int_i0_i27.GSR = "DISABLED";
    FD1P3AX A_int_i0_i26 (.D(alu_a[26]), .SP(n73811), .CK(clock), .Q(A_int[26]));
    defparam A_int_i0_i26.GSR = "DISABLED";
    FD1P3AX A_int_i0_i25 (.D(alu_a[25]), .SP(n73811), .CK(clock), .Q(A_int[25]));
    defparam A_int_i0_i25.GSR = "DISABLED";
    FD1P3AX A_int_i0_i24 (.D(alu_a[24]), .SP(n73811), .CK(clock), .Q(A_int[24]));
    defparam A_int_i0_i24.GSR = "DISABLED";
    FD1P3AX A_int_i0_i23 (.D(alu_a[23]), .SP(n73811), .CK(clock), .Q(A_int[23]));
    defparam A_int_i0_i23.GSR = "DISABLED";
    FD1P3AX A_int_i0_i22 (.D(alu_a[22]), .SP(n73811), .CK(clock), .Q(A_int[22]));
    defparam A_int_i0_i22.GSR = "DISABLED";
    FD1P3AX A_int_i0_i21 (.D(alu_a[21]), .SP(n73811), .CK(clock), .Q(A_int[21]));
    defparam A_int_i0_i21.GSR = "DISABLED";
    FD1P3AX A_int_i0_i20 (.D(alu_a[20]), .SP(n73811), .CK(clock), .Q(A_int[20]));
    defparam A_int_i0_i20.GSR = "DISABLED";
    FD1P3AX A_int_i0_i19 (.D(alu_a[19]), .SP(n73811), .CK(clock), .Q(A_int[19]));
    defparam A_int_i0_i19.GSR = "DISABLED";
    FD1P3AX A_int_i0_i18 (.D(alu_a[18]), .SP(n73811), .CK(clock), .Q(A_int[18]));
    defparam A_int_i0_i18.GSR = "DISABLED";
    FD1P3AX A_int_i0_i17 (.D(alu_a[17]), .SP(n73811), .CK(clock), .Q(A_int[17]));
    defparam A_int_i0_i17.GSR = "DISABLED";
    FD1P3AX A_int_i0_i16 (.D(alu_a[16]), .SP(n73811), .CK(clock), .Q(A_int[16]));
    defparam A_int_i0_i16.GSR = "DISABLED";
    FD1P3AX A_int_i0_i15 (.D(alu_a[15]), .SP(n73811), .CK(clock), .Q(A_int[15]));
    defparam A_int_i0_i15.GSR = "DISABLED";
    FD1P3AX A_int_i0_i14 (.D(alu_a[14]), .SP(n73811), .CK(clock), .Q(A_int[14]));
    defparam A_int_i0_i14.GSR = "DISABLED";
    FD1P3AX A_int_i0_i13 (.D(alu_a[13]), .SP(n73811), .CK(clock), .Q(A_int[13]));
    defparam A_int_i0_i13.GSR = "DISABLED";
    FD1P3AX A_int_i0_i12 (.D(alu_a[12]), .SP(n73811), .CK(clock), .Q(\A_int[12] ));
    defparam A_int_i0_i12.GSR = "DISABLED";
    FD1P3AX A_int_i0_i11 (.D(alu_a[11]), .SP(n73811), .CK(clock), .Q(\A_int[11] ));
    defparam A_int_i0_i11.GSR = "DISABLED";
    FD1P3AX A_int_i0_i10 (.D(alu_a[10]), .SP(n73811), .CK(clock), .Q(\A_int[10] ));
    defparam A_int_i0_i10.GSR = "DISABLED";
    FD1P3AX A_int_i0_i9 (.D(alu_a[9]), .SP(n73811), .CK(clock), .Q(A_int[9]));
    defparam A_int_i0_i9.GSR = "DISABLED";
    FD1P3AX A_int_i0_i8 (.D(alu_a[8]), .SP(n73811), .CK(clock), .Q(A_int[8]));
    defparam A_int_i0_i8.GSR = "DISABLED";
    FD1P3AX A_int_i0_i7 (.D(alu_a[7]), .SP(n73811), .CK(clock), .Q(A_int[7]));
    defparam A_int_i0_i7.GSR = "DISABLED";
    FD1P3AX A_int_i0_i6 (.D(alu_a[6]), .SP(n73811), .CK(clock), .Q(A_int[6]));
    defparam A_int_i0_i6.GSR = "DISABLED";
    FD1P3AX A_int_i0_i5 (.D(alu_a[5]), .SP(n73811), .CK(clock), .Q(A_int[5]));
    defparam A_int_i0_i5.GSR = "DISABLED";
    FD1P3AX A_int_i0_i4 (.D(alu_a[4]), .SP(n73811), .CK(clock), .Q(A_int[4]));
    defparam A_int_i0_i4.GSR = "DISABLED";
    FD1P3AX A_int_i0_i3 (.D(alu_a[3]), .SP(n73811), .CK(clock), .Q(A_int[3]));
    defparam A_int_i0_i3.GSR = "DISABLED";
    FD1P3AX A_int_i0_i2 (.D(alu_a[2]), .SP(n73811), .CK(clock), .Q(A_int[2]));
    defparam A_int_i0_i2.GSR = "DISABLED";
    FD1P3AX A_int_i0_i1 (.D(alu_a[1]), .SP(n73811), .CK(clock), .Q(A_int[1]));
    defparam A_int_i0_i1.GSR = "DISABLED";
    FD1P3AX FP_Z_i0_i31 (.D(sign), .SP(n73811), .CK(clock), .Q(sub_c[31]));
    defparam FP_Z_i0_i31.GSR = "DISABLED";
    FD1P3AX B_int_i0_i31 (.D(alu_b[31]), .SP(sub_ce), .CK(clock), .Q(B_int[31]));
    defparam B_int_i0_i31.GSR = "DISABLED";
    FD1P3AX B_int_i0_i30 (.D(alu_b[30]), .SP(sub_ce), .CK(clock), .Q(B_int[30]));
    defparam B_int_i0_i30.GSR = "DISABLED";
    FD1P3AX B_int_i0_i29 (.D(alu_b[29]), .SP(sub_ce), .CK(clock), .Q(B_int[29]));
    defparam B_int_i0_i29.GSR = "DISABLED";
    FD1P3AX B_int_i0_i28 (.D(alu_b[28]), .SP(sub_ce), .CK(clock), .Q(B_int[28]));
    defparam B_int_i0_i28.GSR = "DISABLED";
    FD1P3AX B_int_i0_i27 (.D(alu_b[27]), .SP(sub_ce), .CK(clock), .Q(B_int[27]));
    defparam B_int_i0_i27.GSR = "DISABLED";
    FD1P3AX B_int_i0_i26 (.D(alu_b[26]), .SP(sub_ce), .CK(clock), .Q(B_int[26]));
    defparam B_int_i0_i26.GSR = "DISABLED";
    FD1P3AX B_int_i0_i25 (.D(alu_b[25]), .SP(sub_ce), .CK(clock), .Q(B_int[25]));
    defparam B_int_i0_i25.GSR = "DISABLED";
    FD1P3AX B_int_i0_i24 (.D(alu_b[24]), .SP(sub_ce), .CK(clock), .Q(B_int[24]));
    defparam B_int_i0_i24.GSR = "DISABLED";
    FD1P3AX B_int_i0_i23 (.D(alu_b[23]), .SP(sub_ce), .CK(clock), .Q(B_int[23]));
    defparam B_int_i0_i23.GSR = "DISABLED";
    FD1P3AX B_int_i0_i22 (.D(alu_b[22]), .SP(sub_ce), .CK(clock), .Q(B_int[22]));
    defparam B_int_i0_i22.GSR = "DISABLED";
    FD1P3AX B_int_i0_i21 (.D(alu_b[21]), .SP(sub_ce), .CK(clock), .Q(B_int[21]));
    defparam B_int_i0_i21.GSR = "DISABLED";
    FD1P3AX B_int_i0_i20 (.D(alu_b[20]), .SP(sub_ce), .CK(clock), .Q(B_int[20]));
    defparam B_int_i0_i20.GSR = "DISABLED";
    FD1P3AX B_int_i0_i19 (.D(alu_b[19]), .SP(sub_ce), .CK(clock), .Q(B_int[19]));
    defparam B_int_i0_i19.GSR = "DISABLED";
    FD1P3AX B_int_i0_i18 (.D(alu_b[18]), .SP(sub_ce), .CK(clock), .Q(B_int[18]));
    defparam B_int_i0_i18.GSR = "DISABLED";
    FD1P3AX B_int_i0_i17 (.D(alu_b[17]), .SP(sub_ce), .CK(clock), .Q(B_int[17]));
    defparam B_int_i0_i17.GSR = "DISABLED";
    FD1P3AX B_int_i0_i16 (.D(alu_b[16]), .SP(sub_ce), .CK(clock), .Q(B_int[16]));
    defparam B_int_i0_i16.GSR = "DISABLED";
    FD1P3AX B_int_i0_i15 (.D(alu_b[15]), .SP(sub_ce), .CK(clock), .Q(B_int[15]));
    defparam B_int_i0_i15.GSR = "DISABLED";
    FD1P3AX B_int_i0_i14 (.D(alu_b[14]), .SP(sub_ce), .CK(clock), .Q(B_int[14]));
    defparam B_int_i0_i14.GSR = "DISABLED";
    FD1P3AX B_int_i0_i13 (.D(alu_b[13]), .SP(sub_ce), .CK(clock), .Q(B_int[13]));
    defparam B_int_i0_i13.GSR = "DISABLED";
    FD1P3AX B_int_i0_i12 (.D(alu_b[12]), .SP(sub_ce), .CK(clock), .Q(\B_int[12] ));
    defparam B_int_i0_i12.GSR = "DISABLED";
    FD1P3AX B_int_i0_i11 (.D(alu_b[11]), .SP(sub_ce), .CK(clock), .Q(\B_int[11] ));
    defparam B_int_i0_i11.GSR = "DISABLED";
    FD1P3AX B_int_i0_i10 (.D(alu_b[10]), .SP(sub_ce), .CK(clock), .Q(\B_int[10] ));
    defparam B_int_i0_i10.GSR = "DISABLED";
    FD1P3AX B_int_i0_i9 (.D(alu_b[9]), .SP(sub_ce), .CK(clock), .Q(B_int[9]));
    defparam B_int_i0_i9.GSR = "DISABLED";
    FD1P3AX B_int_i0_i8 (.D(alu_b[8]), .SP(sub_ce), .CK(clock), .Q(B_int[8]));
    defparam B_int_i0_i8.GSR = "DISABLED";
    FD1P3AX B_int_i0_i7 (.D(alu_b[7]), .SP(sub_ce), .CK(clock), .Q(B_int[7]));
    defparam B_int_i0_i7.GSR = "DISABLED";
    FD1P3AX B_int_i0_i6 (.D(alu_b[6]), .SP(sub_ce), .CK(clock), .Q(B_int[6]));
    defparam B_int_i0_i6.GSR = "DISABLED";
    FD1P3AX B_int_i0_i5 (.D(alu_b[5]), .SP(sub_ce), .CK(clock), .Q(B_int[5]));
    defparam B_int_i0_i5.GSR = "DISABLED";
    FD1P3AX B_int_i0_i4 (.D(alu_b[4]), .SP(sub_ce), .CK(clock), .Q(B_int[4]));
    defparam B_int_i0_i4.GSR = "DISABLED";
    FD1P3AX B_int_i0_i3 (.D(alu_b[3]), .SP(sub_ce), .CK(clock), .Q(B_int[3]));
    defparam B_int_i0_i3.GSR = "DISABLED";
    FD1P3AX B_int_i0_i2 (.D(alu_b[2]), .SP(sub_ce), .CK(clock), .Q(B_int[2]));
    defparam B_int_i0_i2.GSR = "DISABLED";
    FD1P3AX B_int_i0_i1 (.D(alu_b[1]), .SP(sub_ce), .CK(clock), .Q(B_int[1]));
    defparam B_int_i0_i1.GSR = "DISABLED";
    LUT4 n70717_bdd_3_lut (.A(n70717), .B(n73142), .C(addSubAB[27]), .Z(frac_add_Norm1[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70717_bdd_3_lut.init = 16'hcaca;
    PFUMX i57283 (.BLUT(n73141), .ALUT(n70717), .C0(n67674), .Z(n73142));
    LUT4 n70717_bdd_3_lut_57285 (.A(n70717), .B(n73140), .C(n61), .Z(n73141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70717_bdd_3_lut_57285.init = 16'hcaca;
    LUT4 i1_4_lut_adj_919 (.A(n41776), .B(n70837), .C(diffExp[4]), .D(n7), 
         .Z(n21699)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_919.init = 16'hccc6;
    CCU2D sub_214_add_2_21 (.A0(B_int[19]), .B0(A_int[19]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[20]), .B1(A_int[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61564), .COUT(n61565), .S0(subBAExpEq[22]), 
          .S1(subBAExpEq[23]));
    defparam sub_214_add_2_21.INIT0 = 16'h5999;
    defparam sub_214_add_2_21.INIT1 = 16'h5999;
    defparam sub_214_add_2_21.INJECT1_0 = "NO";
    defparam sub_214_add_2_21.INJECT1_1 = "NO";
    PFUMX i57281 (.BLUT(n451[3]), .ALUT(n73139), .C0(n448), .Z(n73140));
    LUT4 i1_2_lut_rep_706_3_lut_4_lut (.A(n61), .B(n67674), .C(addSubAB[27]), 
         .D(n70738), .Z(n70676)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_706_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_751_2_lut_3_lut (.A(n61), .B(n67674), .C(n70738), 
         .Z(n70721)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_751_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_739_3_lut_3_lut_4_lut (.A(n61), .B(n67674), .C(n70738), 
         .D(addSubAB[0]), .Z(n70709)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_739_3_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_adj_920 (.A(n70763), .B(n70837), .C(n41584), .D(n7), 
         .Z(n21717)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_920.init = 16'hcc9c;
    LUT4 i1_2_lut_rep_747_3_lut_3_lut_4_lut (.A(n61), .B(n67674), .C(n70738), 
         .D(addSubAB[2]), .Z(n70717)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_747_3_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i29933_2_lut_rep_748_3_lut_3_lut_4_lut (.A(n61), .B(n67674), .C(n70738), 
         .D(addSubAB[1]), .Z(n70718)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i29933_2_lut_rep_748_3_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 n476_bdd_4_lut (.A(n451[3]), .B(n70717), .C(subBAExpEq[27]), 
         .D(n70837), .Z(n73139)) /* synthesis lut_function=(A (B+(C+(D)))+!A !((C+(D))+!B)) */ ;
    defparam n476_bdd_4_lut.init = 16'haaac;
    LUT4 i1_4_lut_adj_921 (.A(n15), .B(n70837), .C(n7), .D(n70734), 
         .Z(n21719)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_921.init = 16'hccc6;
    LUT4 i55058_2_lut_rep_759 (.A(n61), .B(n67674), .Z(n70729)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i55058_2_lut_rep_759.init = 16'hdddd;
    LUT4 i1_4_lut_adj_922 (.A(n7), .B(n70837), .C(n66912), .D(diffExp[2]), 
         .Z(n21725)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_922.init = 16'hcc9c;
    LUT4 i1_4_lut_adj_923 (.A(n7), .B(n70837), .C(n66898), .D(diffExp[1]), 
         .Z(n21715)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_923.init = 16'hcc9c;
    LUT4 i2_2_lut_rep_647_3_lut_4_lut_4_lut (.A(n70729), .B(n70634), .C(n73796), 
         .D(n70738), .Z(n70617)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i2_2_lut_rep_647_3_lut_4_lut_4_lut.init = 16'hfbff;
    LUT4 i55057_1_lut_4_lut (.A(n66185), .B(n9_adj_498), .C(n14), .D(n10), 
         .Z(n67674)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i55057_1_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_rep_757 (.A(n66185), .B(n9_adj_498), .C(n14), .D(n10), 
         .Z(n70727)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_rep_757.init = 16'hfffe;
    CCU2D sub_214_add_2_19 (.A0(B_int[17]), .B0(A_int[17]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[18]), .B1(A_int[18]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61563), .COUT(n61564), .S0(subBAExpEq[20]), 
          .S1(subBAExpEq[21]));
    defparam sub_214_add_2_19.INIT0 = 16'h5999;
    defparam sub_214_add_2_19.INIT1 = 16'h5999;
    defparam sub_214_add_2_19.INJECT1_0 = "NO";
    defparam sub_214_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_17 (.A0(B_int[15]), .B0(A_int[15]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[16]), .B1(A_int[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61562), .COUT(n61563), .S0(subBAExpEq[18]), 
          .S1(subBAExpEq[19]));
    defparam sub_214_add_2_17.INIT0 = 16'h5999;
    defparam sub_214_add_2_17.INIT1 = 16'h5999;
    defparam sub_214_add_2_17.INJECT1_0 = "NO";
    defparam sub_214_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_15 (.A0(B_int[13]), .B0(A_int[13]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[14]), .B1(A_int[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61561), .COUT(n61562), .S0(subBAExpEq[16]), 
          .S1(subBAExpEq[17]));
    defparam sub_214_add_2_15.INIT0 = 16'h5999;
    defparam sub_214_add_2_15.INIT1 = 16'h5999;
    defparam sub_214_add_2_15.INJECT1_0 = "NO";
    defparam sub_214_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_13 (.A0(\B_int[11] ), .B0(\A_int[11] ), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\A_int[12] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61560), .COUT(n61561), .S0(subBAExpEq[14]), 
          .S1(subBAExpEq[15]));
    defparam sub_214_add_2_13.INIT0 = 16'h5999;
    defparam sub_214_add_2_13.INIT1 = 16'h5999;
    defparam sub_214_add_2_13.INJECT1_0 = "NO";
    defparam sub_214_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_11 (.A0(B_int[9]), .B0(A_int[9]), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\A_int[10] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61559), .COUT(n61560), .S0(subBAExpEq[12]), 
          .S1(subBAExpEq[13]));
    defparam sub_214_add_2_11.INIT0 = 16'h5999;
    defparam sub_214_add_2_11.INIT1 = 16'h5999;
    defparam sub_214_add_2_11.INJECT1_0 = "NO";
    defparam sub_214_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_9 (.A0(B_int[7]), .B0(A_int[7]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[8]), .B1(A_int[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61558), .COUT(n61559), .S0(subBAExpEq[10]), 
          .S1(subBAExpEq[11]));
    defparam sub_214_add_2_9.INIT0 = 16'h5999;
    defparam sub_214_add_2_9.INIT1 = 16'h5999;
    defparam sub_214_add_2_9.INJECT1_0 = "NO";
    defparam sub_214_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_7 (.A0(B_int[5]), .B0(A_int[5]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[6]), .B1(A_int[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61557), .COUT(n61558), .S0(subBAExpEq[8]), 
          .S1(subBAExpEq[9]));
    defparam sub_214_add_2_7.INIT0 = 16'h5999;
    defparam sub_214_add_2_7.INIT1 = 16'h5999;
    defparam sub_214_add_2_7.INJECT1_0 = "NO";
    defparam sub_214_add_2_7.INJECT1_1 = "NO";
    LUT4 mux_33_i18_3_lut_4_lut (.A(addSubAB[1]), .B(n70721), .C(n70634), 
         .D(n70689), .Z(n243[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_33_i18_3_lut_4_lut.init = 16'hf808;
    CCU2D sub_214_add_2_5 (.A0(B_int[3]), .B0(A_int[3]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[4]), .B1(A_int[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61556), .COUT(n61557), .S0(subBAExpEq[6]), 
          .S1(subBAExpEq[7]));
    defparam sub_214_add_2_5.INIT0 = 16'h5999;
    defparam sub_214_add_2_5.INIT1 = 16'h5999;
    defparam sub_214_add_2_5.INJECT1_0 = "NO";
    defparam sub_214_add_2_5.INJECT1_1 = "NO";
    LUT4 mux_3772_i8_4_lut (.A(frac_Norm2[7]), .B(frac[10]), .C(n70729), 
         .D(n70612), .Z(n10672[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i8_4_lut.init = 16'hcac0;
    LUT4 i7726_3_lut_rep_656_4_lut (.A(addSubAB[1]), .B(n70721), .C(n73796), 
         .D(frac[9]), .Z(n70626)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i7726_3_lut_rep_656_4_lut.init = 16'h8f80;
    LUT4 i7702_3_lut_4_lut (.A(addSubAB[2]), .B(n70721), .C(leadZerosBin[2]), 
         .D(frac[6]), .Z(n66825)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i7702_3_lut_4_lut.init = 16'h8f80;
    LUT4 i7724_3_lut_rep_655_4_lut (.A(addSubAB[2]), .B(n70721), .C(n73796), 
         .D(frac[10]), .Z(n70625)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i7724_3_lut_rep_655_4_lut.init = 16'h8f80;
    LUT4 mux_33_i19_3_lut_4_lut (.A(addSubAB[2]), .B(n70721), .C(n70634), 
         .D(frac[18]), .Z(n243[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_33_i19_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_3772_i7_4_lut (.A(frac_Norm2[6]), .B(frac[9]), .C(n70729), 
         .D(n70612), .Z(n10672[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i7_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i6_4_lut (.A(frac_Norm2[5]), .B(n70698), .C(n70729), 
         .D(n70612), .Z(n10672[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i6_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i5_4_lut (.A(frac_Norm2[4]), .B(n73799), .C(n70729), 
         .D(n70612), .Z(n10672[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i5_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_rep_740 (.A(addSubAB[1]), .B(addSubAB[0]), .Z(n70710)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_740.init = 16'heeee;
    LUT4 mux_33_i17_3_lut_4_lut (.A(addSubAB[0]), .B(n70721), .C(n70634), 
         .D(frac[16]), .Z(n243[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_33_i17_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_31_i9_3_lut_4_lut (.A(addSubAB[0]), .B(n70721), .C(n73796), 
         .D(n70698), .Z(n41732)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_31_i9_3_lut_4_lut.init = 16'h8f80;
    CCU2D add_3121_29 (.A0(A_int[31]), .B0(B_int[31]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61839), 
          .S0(addSubAB[27]));
    defparam add_3121_29.INIT0 = 16'h6999;
    defparam add_3121_29.INIT1 = 16'h0000;
    defparam add_3121_29.INJECT1_0 = "NO";
    defparam add_3121_29.INJECT1_1 = "NO";
    CCU2D add_3121_27 (.A0(n21715), .B0(A_int[22]), .C0(B_int[22]), .D0(diffExpAB[8]), 
          .A1(n70837), .B1(n66221), .C1(GND_net), .D1(GND_net), .CIN(n61838), 
          .COUT(n61839), .S0(addSubAB[25]), .S1(addSubAB[26]));
    defparam add_3121_27.INIT0 = 16'ha599;
    defparam add_3121_27.INIT1 = 16'h9999;
    defparam add_3121_27.INJECT1_0 = "NO";
    defparam add_3121_27.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_3 (.A0(B_int[1]), .B0(A_int[1]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[2]), .B1(A_int[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61555), .COUT(n61556), .S0(subBAExpEq[4]), 
          .S1(subBAExpEq[5]));
    defparam sub_214_add_2_3.INIT0 = 16'h5999;
    defparam sub_214_add_2_3.INIT1 = 16'h5999;
    defparam sub_214_add_2_3.INJECT1_0 = "NO";
    defparam sub_214_add_2_3.INJECT1_1 = "NO";
    LUT4 mux_3772_i4_4_lut (.A(frac_Norm2[3]), .B(frac[6]), .C(n70729), 
         .D(n70612), .Z(n10672[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i4_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i3_4_lut (.A(frac_Norm2[2]), .B(n70699), .C(n70729), 
         .D(n70612), .Z(n10672[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i3_4_lut.init = 16'hcac0;
    LUT4 mux_3772_i2_4_lut (.A(frac_Norm2[1]), .B(n70704), .C(n70729), 
         .D(n70612), .Z(n10672[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3772_i2_4_lut.init = 16'hcac0;
    LUT4 i12429_3_lut (.A(n73810), .B(n731), .C(n66231), .Z(n24092)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i12429_3_lut.init = 16'ha8a8;
    CCU2D add_3121_25 (.A0(n21725), .B0(A_int[20]), .C0(B_int[20]), .D0(diffExpAB[8]), 
          .A1(n21719), .B1(A_int[21]), .C1(B_int[21]), .D1(diffExpAB[8]), 
          .CIN(n61837), .COUT(n61838), .S0(addSubAB[23]), .S1(addSubAB[24]));
    defparam add_3121_25.INIT0 = 16'ha599;
    defparam add_3121_25.INIT1 = 16'ha599;
    defparam add_3121_25.INJECT1_0 = "NO";
    defparam add_3121_25.INJECT1_1 = "NO";
    CCU2D add_3121_23 (.A0(n21739), .B0(diffExpAB[8]), .C0(B_int[18]), 
          .D0(A_int[18]), .A1(n21737), .B1(A_int[19]), .C1(B_int[19]), 
          .D1(diffExpAB[8]), .CIN(n61836), .COUT(n61837), .S0(addSubAB[21]), 
          .S1(addSubAB[22]));
    defparam add_3121_23.INIT0 = 16'ha695;
    defparam add_3121_23.INIT1 = 16'ha599;
    defparam add_3121_23.INJECT1_0 = "NO";
    defparam add_3121_23.INJECT1_1 = "NO";
    CCU2D add_3121_21 (.A0(n21717), .B0(A_int[16]), .C0(B_int[16]), .D0(diffExpAB[8]), 
          .A1(n21727), .B1(A_int[17]), .C1(B_int[17]), .D1(diffExpAB[8]), 
          .CIN(n61835), .COUT(n61836), .S0(addSubAB[19]), .S1(addSubAB[20]));
    defparam add_3121_21.INIT0 = 16'ha599;
    defparam add_3121_21.INIT1 = 16'ha599;
    defparam add_3121_21.INJECT1_0 = "NO";
    defparam add_3121_21.INJECT1_1 = "NO";
    CCU2D add_3121_19 (.A0(n21735), .B0(diffExpAB[8]), .C0(B_int[14]), 
          .D0(A_int[14]), .A1(n21733), .B1(A_int[15]), .C1(B_int[15]), 
          .D1(diffExpAB[8]), .CIN(n61834), .COUT(n61835), .S0(addSubAB[17]), 
          .S1(addSubAB[18]));
    defparam add_3121_19.INIT0 = 16'ha695;
    defparam add_3121_19.INIT1 = 16'ha599;
    defparam add_3121_19.INJECT1_0 = "NO";
    defparam add_3121_19.INJECT1_1 = "NO";
    CCU2D add_3121_17 (.A0(n21743), .B0(diffExpAB[8]), .C0(\B_int[12] ), 
          .D0(\A_int[12] ), .A1(n21729), .B1(A_int[13]), .C1(diffExpAB[8]), 
          .D1(B_int[13]), .CIN(n61833), .COUT(n61834), .S0(addSubAB[15]), 
          .S1(addSubAB[16]));
    defparam add_3121_17.INIT0 = 16'ha695;
    defparam add_3121_17.INIT1 = 16'ha959;
    defparam add_3121_17.INJECT1_0 = "NO";
    defparam add_3121_17.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_924 (.A(addSubAB[2]), .B(n70710), .C(n70721), 
         .D(n70635), .Z(n53)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i2_3_lut_4_lut_adj_924.init = 16'hffe0;
    CCU2D add_3121_15 (.A0(n21723), .B0(\A_int[10] ), .C0(diffExpAB[8]), 
          .D0(\B_int[10] ), .A1(n21721), .B1(diffExpAB[8]), .C1(\B_int[11] ), 
          .D1(\A_int[11] ), .CIN(n61832), .COUT(n61833), .S0(addSubAB[13]), 
          .S1(addSubAB[14]));
    defparam add_3121_15.INIT0 = 16'ha959;
    defparam add_3121_15.INIT1 = 16'ha695;
    defparam add_3121_15.INJECT1_0 = "NO";
    defparam add_3121_15.INJECT1_1 = "NO";
    LUT4 i28078_4_lut_3_lut_4_lut (.A(A_int[31]), .B(B_int[31]), .C(addSubAB[27]), 
         .D(diffExpAB[8]), .Z(sign)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+!(C+(D))))) */ ;
    defparam i28078_4_lut_3_lut_4_lut.init = 16'h333a;
    CCU2D sub_214_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(B_int[0]), .B1(A_int[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61555), .S1(subBAExpEq[3]));
    defparam sub_214_add_2_1.INIT0 = 16'h0000;
    defparam sub_214_add_2_1.INIT1 = 16'h5999;
    defparam sub_214_add_2_1.INJECT1_0 = "NO";
    defparam sub_214_add_2_1.INJECT1_1 = "NO";
    CCU2D add_3121_13 (.A0(n21699), .B0(A_int[8]), .C0(B_int[8]), .D0(diffExpAB[8]), 
          .A1(n21741), .B1(A_int[9]), .C1(B_int[9]), .D1(diffExpAB[8]), 
          .CIN(n61831), .COUT(n61832), .S0(addSubAB[11]), .S1(addSubAB[12]));
    defparam add_3121_13.INIT0 = 16'ha599;
    defparam add_3121_13.INIT1 = 16'ha599;
    defparam add_3121_13.INJECT1_0 = "NO";
    defparam add_3121_13.INJECT1_1 = "NO";
    CCU2D add_3121_11 (.A0(n15599), .B0(A_int[6]), .C0(B_int[6]), .D0(diffExpAB[8]), 
          .A1(n21697), .B1(A_int[7]), .C1(B_int[7]), .D1(diffExpAB[8]), 
          .CIN(n61830), .COUT(n61831), .S0(addSubAB[9]), .S1(addSubAB[10]));
    defparam add_3121_11.INIT0 = 16'ha599;
    defparam add_3121_11.INIT1 = 16'ha599;
    defparam add_3121_11.INJECT1_0 = "NO";
    defparam add_3121_11.INJECT1_1 = "NO";
    CCU2D add_3121_9 (.A0(n21673), .B0(A_int[4]), .C0(B_int[4]), .D0(diffExpAB[8]), 
          .A1(n21731), .B1(A_int[5]), .C1(B_int[5]), .D1(diffExpAB[8]), 
          .CIN(n61829), .COUT(n61830), .S0(addSubAB[7]), .S1(addSubAB[8]));
    defparam add_3121_9.INIT0 = 16'ha599;
    defparam add_3121_9.INIT1 = 16'ha599;
    defparam add_3121_9.INJECT1_0 = "NO";
    defparam add_3121_9.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_9 (.A0(A_int[30]), .B0(B_int[30]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61553), .S0(diffExpAB_c[7]), .S1(diffExpAB[8]));
    defparam sub_210_add_2_9.INIT0 = 16'h5999;
    defparam sub_210_add_2_9.INIT1 = 16'hffff;
    defparam sub_210_add_2_9.INJECT1_0 = "NO";
    defparam sub_210_add_2_9.INJECT1_1 = "NO";
    CCU2D add_3121_7 (.A0(n15583), .B0(A_int[2]), .C0(B_int[2]), .D0(diffExpAB[8]), 
          .A1(n21701), .B1(A_int[3]), .C1(B_int[3]), .D1(diffExpAB[8]), 
          .CIN(n61828), .COUT(n61829), .S0(addSubAB[5]), .S1(addSubAB[6]));
    defparam add_3121_7.INIT0 = 16'ha599;
    defparam add_3121_7.INIT1 = 16'ha599;
    defparam add_3121_7.INJECT1_0 = "NO";
    defparam add_3121_7.INJECT1_1 = "NO";
    CCU2D add_3121_5 (.A0(n21703), .B0(A_int[0]), .C0(B_int[0]), .D0(diffExpAB[8]), 
          .A1(n21707), .B1(A_int[1]), .C1(B_int[1]), .D1(diffExpAB[8]), 
          .CIN(n61827), .COUT(n61828), .S0(addSubAB[3]), .S1(addSubAB[4]));
    defparam add_3121_5.INIT0 = 16'ha599;
    defparam add_3121_5.INIT1 = 16'ha599;
    defparam add_3121_5.INJECT1_0 = "NO";
    defparam add_3121_5.INJECT1_1 = "NO";
    CCU2D add_3121_3 (.A0(efectFracB_align[1]), .B0(n70837), .C0(GND_net), 
          .D0(GND_net), .A1(efectFracB_align[2]), .B1(n70837), .C1(GND_net), 
          .D1(GND_net), .CIN(n61826), .COUT(n61827), .S0(addSubAB[1]), 
          .S1(addSubAB[2]));
    defparam add_3121_3.INIT0 = 16'h6999;
    defparam add_3121_3.INIT1 = 16'h6999;
    defparam add_3121_3.INJECT1_0 = "NO";
    defparam add_3121_3.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_7 (.A0(A_int[28]), .B0(B_int[28]), .C0(GND_net), 
          .D0(GND_net), .A1(A_int[29]), .B1(B_int[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61552), .COUT(n61553), .S0(diffExpAB_c[5]), 
          .S1(diffExpAB_c[6]));
    defparam sub_210_add_2_7.INIT0 = 16'h5999;
    defparam sub_210_add_2_7.INIT1 = 16'h5999;
    defparam sub_210_add_2_7.INJECT1_0 = "NO";
    defparam sub_210_add_2_7.INJECT1_1 = "NO";
    CCU2D add_3121_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(isSUB), .B1(n7), .C1(fracAlign_int[0]), .D1(n70837), .COUT(n61826), 
          .S1(addSubAB[0]));
    defparam add_3121_1.INIT0 = 16'hF000;
    defparam add_3121_1.INIT1 = 16'h56a9;
    defparam add_3121_1.INJECT1_0 = "NO";
    defparam add_3121_1.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_5 (.A0(A_int[26]), .B0(B_int[26]), .C0(GND_net), 
          .D0(GND_net), .A1(A_int[27]), .B1(B_int[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61551), .COUT(n61552), .S0(diffExpAB_c[3]), 
          .S1(diffExpAB_c[4]));
    defparam sub_210_add_2_5.INIT0 = 16'h5999;
    defparam sub_210_add_2_5.INIT1 = 16'h5999;
    defparam sub_210_add_2_5.INJECT1_0 = "NO";
    defparam sub_210_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_3 (.A0(A_int[24]), .B0(B_int[24]), .C0(GND_net), 
          .D0(GND_net), .A1(A_int[25]), .B1(B_int[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61550), .COUT(n61551), .S0(diffExpAB_c[1]), 
          .S1(diffExpAB_c[2]));
    defparam sub_210_add_2_3.INIT0 = 16'h5999;
    defparam sub_210_add_2_3.INIT1 = 16'h5999;
    defparam sub_210_add_2_3.INJECT1_0 = "NO";
    defparam sub_210_add_2_3.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(A_int[27]), .B(A_int[23]), .Z(n10_adj_499)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(A_int[26]), .B(A_int[25]), .C(A_int[28]), .D(A_int[30]), 
         .Z(n14_adj_500)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i7_4_lut_adj_925 (.A(A_int[24]), .B(n14_adj_500), .C(n10_adj_499), 
         .D(A_int[29]), .Z(expA_FF)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_925.init = 16'h8000;
    LUT4 i2_2_lut_adj_926 (.A(B_int[25]), .B(B_int[27]), .Z(n10_adj_501)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_926.init = 16'h8888;
    LUT4 i6_4_lut_adj_927 (.A(B_int[26]), .B(B_int[24]), .C(B_int[28]), 
         .D(B_int[30]), .Z(n14_adj_502)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_927.init = 16'h8000;
    LUT4 i7_4_lut_adj_928 (.A(B_int[23]), .B(n14_adj_502), .C(n10_adj_501), 
         .D(B_int[29]), .Z(expB_FF)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_928.init = 16'h8000;
    LUT4 i18_4_lut (.A(frac[9]), .B(n70677), .C(n73799), .D(\frac[15] ), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(n73798), .B(n44), .C(n34), .D(n70717), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(n70709), .B(n70837), .C(n70688), .D(frac[26]), 
         .Z(n41)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(frac[3]), .B(n70698), .C(n70687), .D(n70689), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(n41), .B(n48), .C(n31), .D(n32), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(n70699), .B(frac[21]), .C(n70680), .D(frac[10]), 
         .Z(n45)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i25_4_lut (.A(n45), .B(n50), .C(n39), .D(n40), .Z(n93)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(n8351[3]), .B(n8351[2]), .Z(n10_adj_503)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i7_4_lut_adj_929 (.A(n8351[1]), .B(n8351[6]), .C(n8351[5]), .D(n10_adj_503), 
         .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_929.init = 16'h8000;
    LUT4 i6_4_lut_adj_930 (.A(n8351[0]), .B(n8351[7]), .C(n8351[4]), .D(n93), 
         .Z(n15_adj_504)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_930.init = 16'h8000;
    LUT4 i2_4_lut (.A(expB_FF), .B(n15_adj_504), .C(expA_FF), .D(n16), 
         .Z(n22573)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_931 (.A(expA_FF), .B(n70837), .C(expB_FF), .D(n22573), 
         .Z(n731)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_931.init = 16'hde5a;
    CCU2D sub_210_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[23]), .B1(B_int[23]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61550), .S1(diffExpAB_c[0]));
    defparam sub_210_add_2_1.INIT0 = 16'h0000;
    defparam sub_210_add_2_1.INIT1 = 16'h5999;
    defparam sub_210_add_2_1.INJECT1_0 = "NO";
    defparam sub_210_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_932 (.A(expB_FF), .B(expA_FF), .C(n66185), .D(n66199), 
         .Z(n4_adj_505)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_932.init = 16'heca0;
    LUT4 i2_4_lut_adj_933 (.A(expB_FF), .B(n4_adj_505), .C(n70837), .D(expA_FF), 
         .Z(n66231)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i2_4_lut_adj_933.init = 16'hcecc;
    LUT4 mux_51_i4_3_lut (.A(addSubAB[3]), .B(subBAExpEq[3]), .C(n70738), 
         .Z(n451[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i4_3_lut.init = 16'hacac;
    LUT4 mux_51_i5_3_lut (.A(addSubAB[4]), .B(subBAExpEq[4]), .C(n70738), 
         .Z(n451[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i5_3_lut.init = 16'hacac;
    LUT4 mux_51_i6_3_lut (.A(addSubAB[5]), .B(subBAExpEq[5]), .C(n70738), 
         .Z(n451[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i6_3_lut.init = 16'hacac;
    LUT4 mux_51_i12_3_lut (.A(addSubAB[11]), .B(subBAExpEq[11]), .C(n70738), 
         .Z(n451[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i12_3_lut.init = 16'hacac;
    LUT4 mux_51_i8_3_lut (.A(addSubAB[7]), .B(subBAExpEq[7]), .C(n70738), 
         .Z(n451[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i8_3_lut.init = 16'hacac;
    CCU2D add_72_23 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[24]), 
          .D0(frac_add_Norm1[24]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[25]), 
          .D1(frac_add_Norm1[25]), .CIN(n61548), .S0(frac_Norm2[21]), 
          .S1(frac_Norm2[22]));
    defparam add_72_23.INIT0 = 16'hf690;
    defparam add_72_23.INIT1 = 16'hf690;
    defparam add_72_23.INJECT1_0 = "NO";
    defparam add_72_23.INJECT1_1 = "NO";
    LUT4 mux_51_i9_3_lut (.A(addSubAB[8]), .B(subBAExpEq[8]), .C(n70738), 
         .Z(n451[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i9_3_lut.init = 16'hacac;
    LUT4 mux_51_i10_3_lut (.A(addSubAB[9]), .B(subBAExpEq[9]), .C(n70738), 
         .Z(n451[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i10_3_lut.init = 16'hacac;
    LUT4 mux_51_i11_3_lut (.A(addSubAB[10]), .B(subBAExpEq[10]), .C(n70738), 
         .Z(n451[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i11_3_lut.init = 16'hacac;
    CCU2D add_72_21 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[22]), 
          .D0(frac_add_Norm1[22]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[23]), 
          .D1(frac_add_Norm1[23]), .CIN(n61547), .COUT(n61548), .S0(frac_Norm2[19]), 
          .S1(frac_Norm2[20]));
    defparam add_72_21.INIT0 = 16'hf690;
    defparam add_72_21.INIT1 = 16'hf690;
    defparam add_72_21.INJECT1_0 = "NO";
    defparam add_72_21.INJECT1_1 = "NO";
    LUT4 mux_51_i22_3_lut (.A(addSubAB[21]), .B(subBAExpEq[21]), .C(n70738), 
         .Z(n451[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i22_3_lut.init = 16'hacac;
    LUT4 mux_51_i23_3_lut (.A(addSubAB[22]), .B(subBAExpEq[22]), .C(n70738), 
         .Z(n451[22])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i23_3_lut.init = 16'hacac;
    LUT4 mux_52_i23_3_lut (.A(A_int[19]), .B(n451[22]), .C(n70727), .Z(n480[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i23_3_lut.init = 16'hcaca;
    LUT4 mux_51_i18_3_lut (.A(addSubAB[17]), .B(subBAExpEq[17]), .C(n70738), 
         .Z(n451[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i18_3_lut.init = 16'hacac;
    LUT4 mux_51_i17_3_lut (.A(addSubAB[16]), .B(subBAExpEq[16]), .C(n70738), 
         .Z(n451[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i17_3_lut.init = 16'hacac;
    LUT4 mux_52_i18_3_lut (.A(A_int[14]), .B(n451[17]), .C(n70727), .Z(n480[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i18_3_lut.init = 16'hcaca;
    CCU2D add_72_19 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[20]), 
          .D0(frac_add_Norm1[20]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[21]), 
          .D1(frac_add_Norm1[21]), .CIN(n61546), .COUT(n61547), .S0(frac_Norm2[17]), 
          .S1(frac_Norm2[18]));
    defparam add_72_19.INIT0 = 16'hf690;
    defparam add_72_19.INIT1 = 16'hf690;
    defparam add_72_19.INJECT1_0 = "NO";
    defparam add_72_19.INJECT1_1 = "NO";
    LUT4 mux_51_i16_3_lut (.A(addSubAB[15]), .B(subBAExpEq[15]), .C(n70738), 
         .Z(n451[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i16_3_lut.init = 16'hacac;
    LUT4 mux_52_i16_3_lut (.A(\A_int[12] ), .B(n451[15]), .C(n70727), 
         .Z(n493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i16_3_lut.init = 16'hcaca;
    LUT4 mux_51_i26_3_lut (.A(addSubAB[25]), .B(subBAExpEq[25]), .C(n70738), 
         .Z(n451[25])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i26_3_lut.init = 16'hacac;
    LUT4 mux_52_i26_3_lut (.A(A_int[22]), .B(n451[25]), .C(n70727), .Z(n480[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i26_3_lut.init = 16'hcaca;
    LUT4 mux_51_i24_3_lut (.A(addSubAB[23]), .B(subBAExpEq[23]), .C(n70738), 
         .Z(n451[23])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i24_3_lut.init = 16'hacac;
    CCU2D add_72_17 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[18]), 
          .D0(frac_add_Norm1[18]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[19]), 
          .D1(frac_add_Norm1[19]), .CIN(n61545), .COUT(n61546), .S0(frac_Norm2[15]), 
          .S1(frac_Norm2[16]));
    defparam add_72_17.INIT0 = 16'hf690;
    defparam add_72_17.INIT1 = 16'hf690;
    defparam add_72_17.INJECT1_0 = "NO";
    defparam add_72_17.INJECT1_1 = "NO";
    LUT4 mux_51_i25_3_lut (.A(addSubAB[24]), .B(subBAExpEq[24]), .C(n70738), 
         .Z(n451[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i25_3_lut.init = 16'hacac;
    LUT4 mux_52_i25_3_lut (.A(A_int[21]), .B(n451[24]), .C(n70727), .Z(n480[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i25_3_lut.init = 16'hcaca;
    LUT4 mux_52_i24_3_lut (.A(A_int[20]), .B(n451[23]), .C(n70727), .Z(n480[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i24_3_lut.init = 16'hcaca;
    LUT4 i13_2_lut_3_lut_4_lut (.A(n70693), .B(n70692), .C(frac[6]), .D(frac[12]), 
         .Z(n39)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i27996_2_lut_rep_677_3_lut_4_lut (.A(n70693), .B(n70692), .C(n22515), 
         .D(n70658), .Z(n70647)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i27996_2_lut_rep_677_3_lut_4_lut.init = 16'hf0e0;
    CCU2D add_72_15 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[16]), 
          .D0(frac_add_Norm1[16]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[17]), 
          .D1(frac_add_Norm1[17]), .CIN(n61544), .COUT(n61545), .S0(frac_Norm2[13]), 
          .S1(frac_Norm2[14]));
    defparam add_72_15.INIT0 = 16'hf690;
    defparam add_72_15.INIT1 = 16'hf690;
    defparam add_72_15.INJECT1_0 = "NO";
    defparam add_72_15.INJECT1_1 = "NO";
    LUT4 mux_51_i13_3_lut (.A(addSubAB[12]), .B(subBAExpEq[12]), .C(n70738), 
         .Z(n451[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i13_3_lut.init = 16'hacac;
    LUT4 mux_51_i15_3_lut (.A(addSubAB[14]), .B(subBAExpEq[14]), .C(n70738), 
         .Z(n451[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i15_3_lut.init = 16'hacac;
    LUT4 mux_51_i14_3_lut (.A(addSubAB[13]), .B(subBAExpEq[13]), .C(n70738), 
         .Z(n466)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i14_3_lut.init = 16'hacac;
    CCU2D add_72_13 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[14]), 
          .D0(frac_add_Norm1[14]), .A1(n41812), .B1(n70634), .C1(frac_add_Norm1[15]), 
          .D1(n70837), .CIN(n61543), .COUT(n61544), .S0(frac_Norm2[11]), 
          .S1(frac_Norm2[12]));
    defparam add_72_13.INIT0 = 16'hf690;
    defparam add_72_13.INIT1 = 16'hf088;
    defparam add_72_13.INJECT1_0 = "NO";
    defparam add_72_13.INJECT1_1 = "NO";
    LUT4 mux_52_i15_3_lut (.A(\A_int[11] ), .B(n451[14]), .C(n70727), 
         .Z(n480[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_720_3_lut (.A(n70693), .B(n70692), .C(frac[12]), 
         .Z(n70690)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_720_3_lut.init = 16'hfefe;
    LUT4 mux_52_i13_3_lut (.A(A_int[9]), .B(n451[12]), .C(n70727), .Z(n480[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i13_3_lut.init = 16'hcaca;
    LUT4 mux_51_i21_3_lut (.A(addSubAB[20]), .B(subBAExpEq[20]), .C(n70738), 
         .Z(n451[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i21_3_lut.init = 16'hacac;
    LUT4 mux_51_i19_3_lut (.A(addSubAB[18]), .B(subBAExpEq[18]), .C(n70738), 
         .Z(n451[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i19_3_lut.init = 16'hacac;
    LUT4 i5_2_lut (.A(A_int[15]), .B(\A_int[12] ), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i15_4_lut_adj_934 (.A(A_int[16]), .B(A_int[21]), .C(A_int[3]), 
         .D(A_int[18]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_934.init = 16'hfffe;
    LUT4 i1_2_lut_adj_935 (.A(A_int[1]), .B(A_int[14]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_935.init = 16'heeee;
    LUT4 i13_4_lut (.A(A_int[0]), .B(\A_int[10] ), .C(A_int[19]), .D(A_int[6]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut_adj_936 (.A(A_int[4]), .B(n38), .C(n28), .D(A_int[22]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_936.init = 16'hfffe;
    CCU2D add_72_11 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[12]), 
          .D0(frac_add_Norm1[12]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[13]), 
          .D1(frac_add_Norm1[13]), .CIN(n61542), .COUT(n61543), .S0(frac_Norm2[9]), 
          .S1(frac_Norm2[10]));
    defparam add_72_11.INIT0 = 16'hf690;
    defparam add_72_11.INIT1 = 16'hf690;
    defparam add_72_11.INJECT1_0 = "NO";
    defparam add_72_11.INJECT1_1 = "NO";
    LUT4 i9_2_lut (.A(A_int[20]), .B(A_int[8]), .Z(n32_adj_506)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(A_int[9]), .B(A_int[2]), .C(A_int[5]), .D(A_int[17]), 
         .Z(n40_adj_507)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(A_int[13]), .B(n42), .C(n36), .D(n24), .Z(n44_adj_508)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(\A_int[11] ), .B(A_int[7]), .Z(n31_adj_509)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i22_4_lut_adj_937 (.A(n31_adj_509), .B(n44_adj_508), .C(n40_adj_507), 
         .D(n32_adj_506), .Z(n66199)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut_adj_937.init = 16'hfffe;
    LUT4 i2_2_lut_adj_938 (.A(A_int[24]), .B(A_int[30]), .Z(n10_adj_510)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_938.init = 16'heeee;
    LUT4 i6_4_lut_adj_939 (.A(A_int[28]), .B(A_int[23]), .C(A_int[26]), 
         .D(A_int[27]), .Z(n14_adj_511)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_939.init = 16'hfffe;
    LUT4 i1_2_lut_adj_940 (.A(A_int[25]), .B(A_int[29]), .Z(n9_adj_512)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_940.init = 16'heeee;
    LUT4 i1_4_lut_adj_941 (.A(n66199), .B(n9_adj_512), .C(n14_adj_511), 
         .D(n10_adj_510), .Z(n61)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_941.init = 16'hfffe;
    LUT4 mux_51_i20_3_lut (.A(addSubAB[19]), .B(subBAExpEq[19]), .C(n70738), 
         .Z(n451[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i20_3_lut.init = 16'hacac;
    LUT4 mux_52_i20_3_lut (.A(A_int[16]), .B(n451[19]), .C(n70727), .Z(n480[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i20_3_lut.init = 16'hcaca;
    LUT4 mux_52_i19_3_lut (.A(A_int[15]), .B(n451[18]), .C(n70727), .Z(n480[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i19_3_lut.init = 16'hcaca;
    LUT4 mux_52_i21_3_lut (.A(A_int[17]), .B(n451[20]), .C(n70727), .Z(n480[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i21_3_lut.init = 16'hcaca;
    LUT4 mux_52_i12_3_lut (.A(A_int[8]), .B(n451[11]), .C(n70727), .Z(n480[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i12_3_lut.init = 16'hcaca;
    LUT4 mux_52_i11_3_lut (.A(A_int[7]), .B(n451[10]), .C(n70727), .Z(n480[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i11_3_lut.init = 16'hcaca;
    LUT4 mux_52_i10_3_lut (.A(A_int[6]), .B(n451[9]), .C(n70727), .Z(n480[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i10_3_lut.init = 16'hcaca;
    LUT4 mux_52_i9_3_lut (.A(A_int[5]), .B(n451[8]), .C(n70727), .Z(n480[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i9_3_lut.init = 16'hcaca;
    CCU2D add_72_9 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[10]), 
          .D0(frac_add_Norm1[10]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[11]), 
          .D1(frac_add_Norm1[11]), .CIN(n61541), .COUT(n61542), .S0(frac_Norm2[7]), 
          .S1(frac_Norm2[8]));
    defparam add_72_9.INIT0 = 16'hf690;
    defparam add_72_9.INIT1 = 16'hf690;
    defparam add_72_9.INJECT1_0 = "NO";
    defparam add_72_9.INJECT1_1 = "NO";
    LUT4 i29849_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[21]), 
         .D(n451[20]), .Z(n41444)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29849_3_lut_4_lut.init = 16'hf780;
    LUT4 i29903_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70683), 
         .D(n451[21]), .Z(n41498)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29903_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_52_i8_3_lut (.A(A_int[4]), .B(n451[7]), .C(n70727), .Z(n480[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i8_3_lut.init = 16'hcaca;
    LUT4 i28407_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[26]), 
         .D(n451[25]), .Z(n40000)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i28407_3_lut_4_lut.init = 16'hf780;
    CCU2D add_72_7 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[8]), 
          .D0(frac_add_Norm1[8]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[9]), 
          .D1(frac_add_Norm1[9]), .CIN(n61540), .COUT(n61541), .S0(frac_Norm2[5]), 
          .S1(frac_Norm2[6]));
    defparam add_72_7.INIT0 = 16'hf690;
    defparam add_72_7.INIT1 = 16'hf690;
    defparam add_72_7.INJECT1_0 = "NO";
    defparam add_72_7.INJECT1_1 = "NO";
    LUT4 i5_2_lut_adj_942 (.A(B_int[9]), .B(B_int[5]), .Z(n28_adj_513)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut_adj_942.init = 16'heeee;
    LUT4 i15_4_lut_adj_943 (.A(B_int[2]), .B(B_int[4]), .C(\B_int[10] ), 
         .D(B_int[22]), .Z(n38_adj_514)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_943.init = 16'hfffe;
    LUT4 i1_2_lut_adj_944 (.A(B_int[18]), .B(B_int[1]), .Z(n24_adj_515)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_944.init = 16'heeee;
    LUT4 i13_4_lut_adj_945 (.A(B_int[3]), .B(B_int[19]), .C(B_int[21]), 
         .D(B_int[20]), .Z(n36_adj_516)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_945.init = 16'hfffe;
    LUT4 i19_4_lut_adj_946 (.A(\B_int[12] ), .B(n38_adj_514), .C(n28_adj_513), 
         .D(B_int[0]), .Z(n42_adj_517)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_946.init = 16'hfffe;
    LUT4 i29772_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70699), 
         .D(n451[4]), .Z(n41365)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29772_3_lut_4_lut.init = 16'hf780;
    LUT4 i29780_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[6]), 
         .D(n451[5]), .Z(n41373)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29780_3_lut_4_lut.init = 16'hf780;
    LUT4 i29788_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n73799), 
         .D(n451[6]), .Z(n41381)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29788_3_lut_4_lut.init = 16'hf780;
    LUT4 i9_2_lut_adj_947 (.A(B_int[16]), .B(B_int[17]), .Z(n32_adj_518)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut_adj_947.init = 16'heeee;
    LUT4 i17_4_lut_adj_948 (.A(B_int[13]), .B(B_int[6]), .C(B_int[7]), 
         .D(B_int[15]), .Z(n40_adj_519)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_948.init = 16'hfffe;
    LUT4 i29790_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70698), 
         .D(n451[7]), .Z(n41383)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29790_3_lut_4_lut.init = 16'hf780;
    LUT4 i21_4_lut_adj_949 (.A(\B_int[11] ), .B(n42_adj_517), .C(n36_adj_516), 
         .D(n24_adj_515), .Z(n44_adj_520)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut_adj_949.init = 16'hfffe;
    LUT4 i8_2_lut_adj_950 (.A(B_int[14]), .B(B_int[8]), .Z(n31_adj_521)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut_adj_950.init = 16'heeee;
    LUT4 i29792_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[9]), 
         .D(n451[8]), .Z(n41385)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29792_3_lut_4_lut.init = 16'hf780;
    LUT4 i22_4_lut_adj_951 (.A(n31_adj_521), .B(n44_adj_520), .C(n40_adj_519), 
         .D(n32_adj_518), .Z(n66185)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut_adj_951.init = 16'hfffe;
    CCU2D add_72_5 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[6]), 
          .D0(frac_add_Norm1[6]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[7]), 
          .D1(frac_add_Norm1[7]), .CIN(n61539), .COUT(n61540), .S0(frac_Norm2[3]), 
          .S1(frac_Norm2[4]));
    defparam add_72_5.INIT0 = 16'hf690;
    defparam add_72_5.INIT1 = 16'hf690;
    defparam add_72_5.INJECT1_0 = "NO";
    defparam add_72_5.INJECT1_1 = "NO";
    LUT4 i2_2_lut_adj_952 (.A(B_int[26]), .B(B_int[23]), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_952.init = 16'heeee;
    LUT4 i6_4_lut_adj_953 (.A(B_int[25]), .B(B_int[24]), .C(B_int[27]), 
         .D(B_int[28]), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_953.init = 16'hfffe;
    LUT4 i29798_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[12]), 
         .D(n451[11]), .Z(n41391)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29798_3_lut_4_lut.init = 16'hf780;
    CCU2D add_72_3 (.A0(B_int[31]), .B0(A_int[31]), .C0(frac_sub_Norm1[4]), 
          .D0(frac_add_Norm1[4]), .A1(B_int[31]), .B1(A_int[31]), .C1(frac_sub_Norm1[5]), 
          .D1(frac_add_Norm1[5]), .CIN(n61538), .COUT(n61539), .S0(frac_Norm2[1]), 
          .S1(frac_Norm2[2]));
    defparam add_72_3.INIT0 = 16'hf690;
    defparam add_72_3.INIT1 = 16'hf690;
    defparam add_72_3.INJECT1_0 = "NO";
    defparam add_72_3.INJECT1_1 = "NO";
    CCU2D add_72_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(frac_Norm1[3]), .B1(n70837), .C1(n79), .D1(n63641), .COUT(n61538), 
          .S1(frac_Norm2[0]));
    defparam add_72_1.INIT0 = 16'hF000;
    defparam add_72_1.INIT1 = 16'h596a;
    defparam add_72_1.INJECT1_0 = "NO";
    defparam add_72_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_954 (.A(B_int[30]), .B(B_int[29]), .Z(n9_adj_498)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_954.init = 16'heeee;
    LUT4 i29800_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70692), 
         .D(n451[12]), .Z(n41393)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29800_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_51_i7_3_lut (.A(addSubAB[6]), .B(subBAExpEq[6]), .C(n70738), 
         .Z(n451[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_51_i7_3_lut.init = 16'hacac;
    LUT4 i29802_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70693), 
         .D(n466), .Z(n41395)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29802_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_52_i7_3_lut (.A(A_int[3]), .B(n451[6]), .C(n70727), .Z(n480[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i7_3_lut.init = 16'hcaca;
    LUT4 i29810_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(\frac[15] ), 
         .D(n451[14]), .Z(n41403)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29810_3_lut_4_lut.init = 16'hf780;
    LUT4 i29812_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[16]), 
         .D(n451[15]), .Z(n41405)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29812_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_52_i6_3_lut (.A(A_int[2]), .B(n451[5]), .C(n70727), .Z(n480[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i6_3_lut.init = 16'hcaca;
    LUT4 i29824_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70689), 
         .D(n451[16]), .Z(n41417)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29824_3_lut_4_lut.init = 16'hf780;
    LUT4 i29905_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70681), 
         .D(n451[22]), .Z(n41500)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29905_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_52_i5_3_lut (.A(A_int[1]), .B(n451[4]), .C(n70727), .Z(n480[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_52_i5_3_lut.init = 16'hcaca;
    LUT4 i29847_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70688), 
         .D(n451[19]), .Z(n41442)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29847_3_lut_4_lut.init = 16'hf780;
    LUT4 i29796_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n73798), 
         .D(n451[10]), .Z(n41389)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29796_3_lut_4_lut.init = 16'hf780;
    LUT4 i29845_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70687), 
         .D(n451[18]), .Z(n41440)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29845_3_lut_4_lut.init = 16'hf780;
    LUT4 i28405_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70677), 
         .D(n451[24]), .Z(n39998)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i28405_3_lut_4_lut.init = 16'hf780;
    LUT4 n6_bdd_3_lut_55877_4_lut (.A(n70738), .B(addSubAB[27]), .C(n451[3]), 
         .D(n70704), .Z(n70132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam n6_bdd_3_lut_55877_4_lut.init = 16'hf870;
    LUT4 i28403_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(n70680), 
         .D(n451[23]), .Z(n39996)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i28403_3_lut_4_lut.init = 16'hf780;
    LUT4 i29826_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[18]), 
         .D(n451[17]), .Z(n41419)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29826_3_lut_4_lut.init = 16'hf780;
    LUT4 i29794_3_lut_4_lut (.A(n70738), .B(addSubAB[27]), .C(frac[10]), 
         .D(n451[9]), .Z(n41387)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i29794_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_955 (.A(n70738), .B(addSubAB[27]), .C(addSubAB[2]), 
         .D(n70710), .Z(n66709)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut_adj_955.init = 16'hff80;
    PFUMX i28360 (.BLUT(n39998), .ALUT(n39999), .C0(n70729), .Z(frac_add_Norm1[24]));
    PFUMX i28362 (.BLUT(n39996), .ALUT(n39997), .C0(n70729), .Z(frac_add_Norm1[23]));
    PFUMX i28364 (.BLUT(n41500), .ALUT(n41501), .C0(n70729), .Z(frac_add_Norm1[22]));
    PFUMX i28370 (.BLUT(n41442), .ALUT(n41443), .C0(n70729), .Z(frac_add_Norm1[19]));
    PFUMX i28372 (.BLUT(n41440), .ALUT(n41441), .C0(n70729), .Z(frac_add_Norm1[18]));
    PFUMX i28374 (.BLUT(n41419), .ALUT(n41420), .C0(n70729), .Z(frac_add_Norm1[17]));
    PFUMX i28376 (.BLUT(n41417), .ALUT(n41418), .C0(n70729), .Z(frac_add_Norm1[16]));
    PFUMX i28378 (.BLUT(n41405), .ALUT(n41406), .C0(n70729), .Z(frac_add_Norm1[15]));
    PFUMX i28380 (.BLUT(n41403), .ALUT(n41404), .C0(n70729), .Z(frac_add_Norm1[14]));
    PFUMX i28382 (.BLUT(n41395), .ALUT(n41396), .C0(n70729), .Z(frac_add_Norm1[13]));
    PFUMX i28384 (.BLUT(n41393), .ALUT(n41394), .C0(n70729), .Z(frac_add_Norm1[12]));
    PFUMX i28386 (.BLUT(n41391), .ALUT(n41392), .C0(n70729), .Z(frac_add_Norm1[11]));
    PFUMX i28388 (.BLUT(n41389), .ALUT(n41390), .C0(n70729), .Z(frac_add_Norm1[10]));
    PFUMX i28390 (.BLUT(n41387), .ALUT(n41388), .C0(n70729), .Z(frac_add_Norm1[9]));
    PFUMX i28392 (.BLUT(n41385), .ALUT(n41386), .C0(n70729), .Z(frac_add_Norm1[8]));
    PFUMX i28394 (.BLUT(n41383), .ALUT(n41384), .C0(n70729), .Z(frac_add_Norm1[7]));
    PFUMX i28396 (.BLUT(n41381), .ALUT(n41382), .C0(n70729), .Z(frac_add_Norm1[6]));
    PFUMX i28398 (.BLUT(n41373), .ALUT(n41374), .C0(n70729), .Z(frac_add_Norm1[5]));
    PFUMX i28400 (.BLUT(n41365), .ALUT(n41366), .C0(n70729), .Z(frac_add_Norm1[4]));
    PFUMX i28358 (.BLUT(n40000), .ALUT(n40001), .C0(n70729), .Z(frac_add_Norm1[25]));
    PFUMX i28366 (.BLUT(n41498), .ALUT(n41499), .C0(n70729), .Z(frac_add_Norm1[21]));
    PFUMX i28368 (.BLUT(n41444), .ALUT(n41445), .C0(n70729), .Z(frac_add_Norm1[20]));
    LUT4 i14_4_lut_adj_956 (.A(n70687), .B(n70677), .C(n70680), .D(frac[6]), 
         .Z(n39_adj_522)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i14_4_lut_adj_956.init = 16'h8000;
    LUT4 i16_4_lut (.A(n70692), .B(frac[18]), .C(n70683), .D(n70681), 
         .Z(n41_adj_523)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut.init = 16'h8000;
    LUT4 i20_4_lut (.A(n39_adj_522), .B(n70689), .C(n30), .D(frac[3]), 
         .Z(n45_adj_524)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20_4_lut.init = 16'h8000;
    LUT4 i19_4_lut_adj_957 (.A(n37), .B(frac[10]), .C(n73799), .D(n70698), 
         .Z(n44_adj_525)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19_4_lut_adj_957.init = 16'h8000;
    LUT4 i23_4_lut (.A(n45_adj_524), .B(n41_adj_523), .C(n33), .D(n34_adj_526), 
         .Z(n48_adj_527)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'h8000;
    LUT4 i18_4_lut_adj_958 (.A(n70717), .B(frac[16]), .C(frac[12]), .D(frac[21]), 
         .Z(n43)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18_4_lut_adj_958.init = 16'h8000;
    LUT4 i63_4_lut (.A(n70676), .B(n43), .C(n48_adj_527), .D(n44_adj_525), 
         .Z(n574)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i63_4_lut.init = 16'heaaa;
    CCU2D sub_211_add_2_9 (.A0(B_int[30]), .B0(A_int[30]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62172), .S0(diffExpBA[7]), .S1(diffExpBA[8]));
    defparam sub_211_add_2_9.INIT0 = 16'h5999;
    defparam sub_211_add_2_9.INIT1 = 16'hffff;
    defparam sub_211_add_2_9.INJECT1_0 = "NO";
    defparam sub_211_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_211_add_2_7 (.A0(B_int[28]), .B0(A_int[28]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[29]), .B1(A_int[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62171), .COUT(n62172), .S0(diffExpBA[5]), 
          .S1(diffExpBA[6]));
    defparam sub_211_add_2_7.INIT0 = 16'h5999;
    defparam sub_211_add_2_7.INIT1 = 16'h5999;
    defparam sub_211_add_2_7.INJECT1_0 = "NO";
    defparam sub_211_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_211_add_2_5 (.A0(B_int[26]), .B0(A_int[26]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[27]), .B1(A_int[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62170), .COUT(n62171), .S0(diffExpBA[3]), 
          .S1(diffExpBA[4]));
    defparam sub_211_add_2_5.INIT0 = 16'h5999;
    defparam sub_211_add_2_5.INIT1 = 16'h5999;
    defparam sub_211_add_2_5.INJECT1_0 = "NO";
    defparam sub_211_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_211_add_2_3 (.A0(B_int[24]), .B0(A_int[24]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[25]), .B1(A_int[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62169), .COUT(n62170), .S0(diffExpBA[1]), 
          .S1(diffExpBA[2]));
    defparam sub_211_add_2_3.INIT0 = 16'h5999;
    defparam sub_211_add_2_3.INIT1 = 16'h5999;
    defparam sub_211_add_2_3.INJECT1_0 = "NO";
    defparam sub_211_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_211_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(B_int[23]), .B1(A_int[23]), .C1(GND_net), .D1(GND_net), 
          .COUT(n62169), .S1(diffExpBA[0]));
    defparam sub_211_add_2_1.INIT0 = 16'h0000;
    defparam sub_211_add_2_1.INIT1 = 16'h5999;
    defparam sub_211_add_2_1.INJECT1_0 = "NO";
    defparam sub_211_add_2_1.INJECT1_1 = "NO";
    CCU2D add_3794_9 (.A0(n70837), .B0(A_int[29]), .C0(B_int[29]), .D0(diffExpAB[8]), 
          .A1(n70837), .B1(A_int[30]), .C1(B_int[30]), .D1(diffExpAB[8]), 
          .CIN(n61621), .S0(n8351[6]), .S1(n8351[7]));
    defparam add_3794_9.INIT0 = 16'ha599;
    defparam add_3794_9.INIT1 = 16'ha599;
    defparam add_3794_9.INJECT1_0 = "NO";
    defparam add_3794_9.INJECT1_1 = "NO";
    CCU2D add_3794_7 (.A0(n41446), .B0(A_int[27]), .C0(B_int[27]), .D0(diffExpAB[8]), 
          .A1(n70837), .B1(A_int[28]), .C1(B_int[28]), .D1(diffExpAB[8]), 
          .CIN(n61620), .COUT(n61621), .S0(n8351[4]), .S1(n8351[5]));
    defparam add_3794_7.INIT0 = 16'ha599;
    defparam add_3794_7.INIT1 = 16'ha599;
    defparam add_3794_7.INJECT1_0 = "NO";
    defparam add_3794_7.INJECT1_1 = "NO";
    CCU2D add_3794_5 (.A0(n41450), .B0(A_int[25]), .C0(B_int[25]), .D0(diffExpAB[8]), 
          .A1(n41448), .B1(A_int[26]), .C1(B_int[26]), .D1(diffExpAB[8]), 
          .CIN(n61619), .COUT(n61620), .S0(n8351[2]), .S1(n8351[3]));
    defparam add_3794_5.INIT0 = 16'ha599;
    defparam add_3794_5.INIT1 = 16'ha599;
    defparam add_3794_5.INJECT1_0 = "NO";
    defparam add_3794_5.INJECT1_1 = "NO";
    CCU2D add_3794_3 (.A0(efectExp[0]), .B0(leadZerosBin[0]), .C0(n574), 
          .D0(n70837), .A1(n41452), .B1(A_int[24]), .C1(B_int[24]), 
          .D1(diffExpAB[8]), .CIN(n61618), .COUT(n61619), .S0(n8351[0]), 
          .S1(n8351[1]));
    defparam add_3794_3.INIT0 = 16'h5a99;
    defparam add_3794_3.INIT1 = 16'ha599;
    defparam add_3794_3.INJECT1_0 = "NO";
    defparam add_3794_3.INJECT1_1 = "NO";
    CCU2D add_3794_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[31]), .B1(B_int[31]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61618));
    defparam add_3794_1.INIT0 = 16'hF000;
    defparam add_3794_1.INIT1 = 16'h6666;
    defparam add_3794_1.INJECT1_0 = "NO";
    defparam add_3794_1.INJECT1_1 = "NO";
    LUT4 i29362_2_lut_3_lut (.A(n70634), .B(n73796), .C(n73799), .Z(n272[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29362_2_lut_3_lut.init = 16'h2020;
    LUT4 i29363_2_lut_3_lut (.A(n70634), .B(n73796), .C(frac[6]), .Z(n272[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29363_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_4_lut_adj_959 (.A(n53), .B(n70837), .C(n62960), .D(n93), 
         .Z(n103)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_959.init = 16'hec00;
    LUT4 i29364_2_lut_3_lut (.A(n70634), .B(n73796), .C(n70699), .Z(n272[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29364_2_lut_3_lut.init = 16'h2020;
    LUT4 i6875_2_lut_3_lut_4_lut (.A(n70634), .B(n73796), .C(leadZerosBin[2]), 
         .D(n70721), .Z(n17520)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i6875_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i29365_2_lut_3_lut (.A(n70634), .B(n73796), .C(n70704), .Z(n272[4])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29365_2_lut_3_lut.init = 16'h2020;
    LUT4 i35_4_lut_4_lut (.A(n330[2]), .B(n18), .C(n66711), .D(leadZerosBin[0]), 
         .Z(n63641)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C (D)))) */ ;
    defparam i35_4_lut_4_lut.init = 16'hc0a8;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut_4_lut (.A(addSubAB[1]), .B(n70721), 
         .C(addSubAB[0]), .D(addSubAB[2]), .Z(n66493)) /* synthesis lut_function=(!(A ((D)+!B)+!A (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h008d;
    \fp_leading_zeros_and_shift(27,8,4)  subtraction_norm (.\A_int[28] (A_int[28]), 
            .\B_int[28] (B_int[28]), .\diffExpAB[8] (diffExpAB[8]), .\efectExp[5] (efectExp[5]), 
            .\A_int[29] (A_int[29]), .\B_int[29] (B_int[29]), .\efectExp[6] (efectExp[6]), 
            .\A_int[30] (A_int[30]), .\B_int[30] (B_int[30]), .\efectExp[7] (efectExp[7]), 
            .n62960(n62960), .\B_int[0] (B_int[0]), .n505(n480[3]), .n61(n61), 
            .\frac[3] (frac[3]), .\frac[21] (frac[21]), .n70699(n70699), 
            .n70634(n70634), .n70688(n70688), .n70704(n70704), .n70687(n70687), 
            .\frac[15] (\frac[15] ), .\leadZerosBin[2] (leadZerosBin[2]), 
            .n70681(n70681), .n73799(n73799), .n70693(n70693), .n70683(n70683), 
            .\frac[6] (frac[6]), .n70717(n70717), .n70635(n70635), .n73796(n73796), 
            .\efectExp[4] (efectExp[4]), .n70782(n70782), .\efectExp[2] (efectExp[2]), 
            .\A_int[27] (A_int[27]), .\B_int[27] (B_int[27]), .\efectExp[0] (efectExp[0]), 
            .\efectExp[1] (efectExp[1]), .\leadZerosBin[1] (leadZerosBin[1]), 
            .\leadZerosBin[0] (leadZerosBin[0]), .\A_int[25] (A_int[25]), 
            .\B_int[25] (B_int[25]), .\A_int[24] (A_int[24]), .\B_int[24] (B_int[24]), 
            .\A_int[23] (A_int[23]), .\B_int[23] (B_int[23]), .n354(n330[4]), 
            .\frac_sub_Norm1[5] (frac_sub_Norm1[5]), .n296(n272[4]), .\addSubAB[0] (addSubAB[0]), 
            .n70617(n70617), .n325(n301[4]), .n66873(n66873), .n4(n4), 
            .n351(n330[7]), .n352(n330[6]), .\frac_sub_Norm1[7] (frac_sub_Norm1[7]), 
            .\frac_sub_Norm1[6] (frac_sub_Norm1[6]), .n66825(n66825), .n323(n301[6]), 
            .n41732(n41732), .n321(n301[8]), .n349(n330[9]), .n70067(n70067), 
            .\A_int[26] (A_int[26]), .\B_int[26] (B_int[26]), .n347(n330[11]), 
            .n41774(n41774), .n345(n330[13]), .n41812(n41812), .\frac_sub_Norm1[14] (frac_sub_Norm1[14]), 
            .n70625(n70625), .n70626(n70626), .\frac_sub_Norm1[17] (frac_sub_Norm1[17]), 
            .\frac_sub_Norm1[16] (frac_sub_Norm1[16]), .\frac[12] (frac[12]), 
            .\frac_sub_Norm1[19] (frac_sub_Norm1[19]), .\frac_sub_Norm1[18] (frac_sub_Norm1[18]), 
            .\frac_sub_Norm1[4] (frac_sub_Norm1[4]), .n70692(n70692), .\frac_sub_Norm1[21] (frac_sub_Norm1[21]), 
            .\frac_sub_Norm1[20] (frac_sub_Norm1[20]), .n255(n243[16]), 
            .n70698(n70698), .\frac_sub_Norm1[23] (frac_sub_Norm1[23]), 
            .\frac_sub_Norm1[22] (frac_sub_Norm1[22]), .n70639(n70639), 
            .n73797(n73797), .n254(n243[17]), .\frac[9] (frac[9]), .\addSubAB[1] (addSubAB[1]), 
            .n70721(n70721), .n70647(n70647), .n53(n53), .n70718(n70718), 
            .n66493(n66493), .\frac_sub_Norm1[24] (frac_sub_Norm1[24]), 
            .n70680(n70680), .\B_int[4] (B_int[4]), .n501(n480[7]), .\B_int[8] (B_int[8]), 
            .n497(n480[11]), .n22515(n22515), .n73798(n73798), .\B_int[1] (B_int[1]), 
            .n504(n480[4]), .n32(n32), .\B_int[2] (B_int[2]), .n503(n480[5]), 
            .\frac[26] (frac[26]), .n30(n30), .\B_int[5] (B_int[5]), .n500(n480[8]), 
            .\addSubAB[26] (addSubAB[26]), .n70729(n70729), .\subBAExpEq[26] (subBAExpEq[26]), 
            .n70738(n70738), .n33(n33), .\B_int[11] (\B_int[11] ), .n494(n480[14]), 
            .n37(n37), .\B_int[9] (B_int[9]), .n496(n480[12]), .\B_int[14] (B_int[14]), 
            .n491(n480[17]), .\frac[16] (frac[16]), .n70689(n70689), .\B_int[17] (B_int[17]), 
            .n488(n480[20]), .n34(n34_adj_526), .\B_int[16] (B_int[16]), 
            .n489(n480[19]), .\frac[18] (frac[18]), .\B_int[15] (B_int[15]), 
            .n490(n480[18]), .\B_int[19] (B_int[19]), .n486(n480[22]), 
            .n34_adj_1(n34), .n70690(n70690), .\B_int[20] (B_int[20]), 
            .n485(n480[23]), .n31(n31), .\B_int[7] (B_int[7]), .n498(n480[10]), 
            .\frac[10] (frac[10]), .\B_int[21] (B_int[21]), .n484(n480[24]), 
            .\B_int[6] (B_int[6]), .n499(n480[9]), .\B_int[3] (B_int[3]), 
            .n502(n480[6]), .n70677(n70677), .\B_int[22] (B_int[22]), 
            .n483(n480[25]), .n253(n243[18]), .n261(n243[10]), .n259(n243[12]), 
            .n258(n243[13]), .n295(n272[5]), .n294(n272[6]), .n319(n301[10]), 
            .n293(n272[7]), .n70658(n70658), .n70691(n70691), .\frac_sub_Norm1[25] (frac_sub_Norm1[25]), 
            .n356(n330[2]), .n70134(n70134), .n70620(n70620), .n70618(n70618));
    \right_shifter(27,8,4)  alignment (.diffExpAB({diffExpAB[8], diffExpAB_c[7:0]}), 
            .diffExpBA({diffExpBA}), .\diffExp[4] (diffExp[4]), .n70763(n70763), 
            .\B_int[21] (B_int[21]), .\A_int[21] (A_int[21]), .\diffExp[1] (diffExp[1]), 
            .\B_int[19] (B_int[19]), .\A_int[19] (A_int[19]), .\B_int[14] (B_int[14]), 
            .\A_int[14] (A_int[14]), .\B_int[15] (B_int[15]), .\A_int[15] (A_int[15]), 
            .\B_int[13] (B_int[13]), .\A_int[13] (A_int[13]), .\B_int[7] (B_int[7]), 
            .\A_int[7] (A_int[7]), .\B_int[4] (B_int[4]), .\A_int[4] (A_int[4]), 
            .\efectFracB[13] (\efectFracB[13] ), .\diffExp[2] (diffExp[2]), 
            .n70734(n70734), .n15(n15), .\efectFracB[15] (\efectFracB[15] ), 
            .\efectFracB[14] (\efectFracB[14] ), .\fracAlign_int[0] (fracAlign_int[0]), 
            .n7(n7), .\efectFracB_align[2] (efectFracB_align[2]), .\efectFracB_align[1] (efectFracB_align[1]), 
            .\B_int[0] (B_int[0]), .\A_int[0] (A_int[0]), .\B_int[1] (B_int[1]), 
            .\A_int[1] (A_int[1]), .\fracAlign_int[4] (fracAlign_int[4]), 
            .\fracAlign_int[3] (fracAlign_int[3]), .\B_int[3] (B_int[3]), 
            .\A_int[3] (A_int[3]), .\B_int[2] (B_int[2]), .\A_int[2] (A_int[2]), 
            .\fracAlign_int[6] (fracAlign_int[6]), .\fracAlign_int[5] (fracAlign_int[5]), 
            .\B_int[5] (B_int[5]), .\A_int[5] (A_int[5]), .\fracAlign_int[8] (fracAlign_int[8]), 
            .\fracAlign_int[7] (fracAlign_int[7]), .\B_int[6] (B_int[6]), 
            .\A_int[6] (A_int[6]), .\fracAlign_int[10] (fracAlign_int[10]), 
            .\fracAlign_int[9] (fracAlign_int[9]), .\B_int[9] (B_int[9]), 
            .\A_int[9] (A_int[9]), .\B_int[8] (B_int[8]), .\A_int[8] (A_int[8]), 
            .\fracAlign_int[12] (fracAlign_int[12]), .n66898(n66898), .n41776(n41776), 
            .\fracAlign_int[14] (fracAlign_int[14]), .\fracAlign_int[13] (fracAlign_int[13]), 
            .\fracAlign_int[16] (fracAlign_int[16]), .\fracAlign_int[15] (fracAlign_int[15]), 
            .\fracAlign_int[18] (fracAlign_int[18]), .\fracAlign_int[17] (fracAlign_int[17]), 
            .\B_int[17] (B_int[17]), .\A_int[17] (A_int[17]), .\B_int[16] (B_int[16]), 
            .\A_int[16] (A_int[16]), .\B_int[18] (B_int[18]), .\A_int[18] (A_int[18]), 
            .\fracAlign_int[20] (fracAlign_int[20]), .n41584(n41584), .\fracAlign_int[22] (fracAlign_int[22]), 
            .\fracAlign_int[21] (fracAlign_int[21]), .\B_int[20] (B_int[20]), 
            .\A_int[20] (A_int[20]), .n66912(n66912), .\B_int[22] (B_int[22]), 
            .\A_int[22] (A_int[22]), .n66221(n66221), .n458(n451[21]), 
            .n70727(n70727), .n61(n61), .\frac[21] (frac[21]), .n463(n451[16]), 
            .\frac[16] (frac[16]));
    
endmodule
//
// Verilog Description of module \fp_leading_zeros_and_shift(27,8,4) 
//

module \fp_leading_zeros_and_shift(27,8,4)  (\A_int[28] , \B_int[28] , \diffExpAB[8] , 
            \efectExp[5] , \A_int[29] , \B_int[29] , \efectExp[6] , 
            \A_int[30] , \B_int[30] , \efectExp[7] , n62960, \B_int[0] , 
            n505, n61, \frac[3] , \frac[21] , n70699, n70634, n70688, 
            n70704, n70687, \frac[15] , \leadZerosBin[2] , n70681, 
            n73799, n70693, n70683, \frac[6] , n70717, n70635, n73796, 
            \efectExp[4] , n70782, \efectExp[2] , \A_int[27] , \B_int[27] , 
            \efectExp[0] , \efectExp[1] , \leadZerosBin[1] , \leadZerosBin[0] , 
            \A_int[25] , \B_int[25] , \A_int[24] , \B_int[24] , \A_int[23] , 
            \B_int[23] , n354, \frac_sub_Norm1[5] , n296, \addSubAB[0] , 
            n70617, n325, n66873, n4, n351, n352, \frac_sub_Norm1[7] , 
            \frac_sub_Norm1[6] , n66825, n323, n41732, n321, n349, 
            n70067, \A_int[26] , \B_int[26] , n347, n41774, n345, 
            n41812, \frac_sub_Norm1[14] , n70625, n70626, \frac_sub_Norm1[17] , 
            \frac_sub_Norm1[16] , \frac[12] , \frac_sub_Norm1[19] , \frac_sub_Norm1[18] , 
            \frac_sub_Norm1[4] , n70692, \frac_sub_Norm1[21] , \frac_sub_Norm1[20] , 
            n255, n70698, \frac_sub_Norm1[23] , \frac_sub_Norm1[22] , 
            n70639, n73797, n254, \frac[9] , \addSubAB[1] , n70721, 
            n70647, n53, n70718, n66493, \frac_sub_Norm1[24] , n70680, 
            \B_int[4] , n501, \B_int[8] , n497, n22515, n73798, 
            \B_int[1] , n504, n32, \B_int[2] , n503, \frac[26] , 
            n30, \B_int[5] , n500, \addSubAB[26] , n70729, \subBAExpEq[26] , 
            n70738, n33, \B_int[11] , n494, n37, \B_int[9] , n496, 
            \B_int[14] , n491, \frac[16] , n70689, \B_int[17] , n488, 
            n34, \B_int[16] , n489, \frac[18] , \B_int[15] , n490, 
            \B_int[19] , n486, n34_adj_1, n70690, \B_int[20] , n485, 
            n31, \B_int[7] , n498, \frac[10] , \B_int[21] , n484, 
            \B_int[6] , n499, \B_int[3] , n502, n70677, \B_int[22] , 
            n483, n253, n261, n259, n258, n295, n294, n319, 
            n293, n70658, n70691, \frac_sub_Norm1[25] , n356, n70134, 
            n70620, n70618);
    input \A_int[28] ;
    input \B_int[28] ;
    input \diffExpAB[8] ;
    output \efectExp[5] ;
    input \A_int[29] ;
    input \B_int[29] ;
    output \efectExp[6] ;
    input \A_int[30] ;
    input \B_int[30] ;
    output \efectExp[7] ;
    output n62960;
    input \B_int[0] ;
    input n505;
    input n61;
    output \frac[3] ;
    input \frac[21] ;
    output n70699;
    output n70634;
    output n70688;
    output n70704;
    output n70687;
    input \frac[15] ;
    output \leadZerosBin[2] ;
    output n70681;
    output n73799;
    output n70693;
    output n70683;
    output \frac[6] ;
    input n70717;
    output n70635;
    output n73796;
    output \efectExp[4] ;
    output n70782;
    output \efectExp[2] ;
    input \A_int[27] ;
    input \B_int[27] ;
    output \efectExp[0] ;
    output \efectExp[1] ;
    output \leadZerosBin[1] ;
    output \leadZerosBin[0] ;
    input \A_int[25] ;
    input \B_int[25] ;
    input \A_int[24] ;
    input \B_int[24] ;
    input \A_int[23] ;
    input \B_int[23] ;
    input n354;
    output \frac_sub_Norm1[5] ;
    input n296;
    input \addSubAB[0] ;
    input n70617;
    output n325;
    output n66873;
    input n4;
    output n351;
    input n352;
    output \frac_sub_Norm1[7] ;
    output \frac_sub_Norm1[6] ;
    input n66825;
    output n323;
    input n41732;
    output n321;
    output n349;
    output n70067;
    input \A_int[26] ;
    input \B_int[26] ;
    output n347;
    output n41774;
    output n345;
    output n41812;
    output \frac_sub_Norm1[14] ;
    input n70625;
    input n70626;
    output \frac_sub_Norm1[17] ;
    output \frac_sub_Norm1[16] ;
    output \frac[12] ;
    output \frac_sub_Norm1[19] ;
    output \frac_sub_Norm1[18] ;
    output \frac_sub_Norm1[4] ;
    input n70692;
    output \frac_sub_Norm1[21] ;
    output \frac_sub_Norm1[20] ;
    input n255;
    output n70698;
    output \frac_sub_Norm1[23] ;
    output \frac_sub_Norm1[22] ;
    output n70639;
    output n73797;
    input n254;
    output \frac[9] ;
    input \addSubAB[1] ;
    input n70721;
    input n70647;
    input n53;
    input n70718;
    input n66493;
    output \frac_sub_Norm1[24] ;
    output n70680;
    input \B_int[4] ;
    input n501;
    input \B_int[8] ;
    input n497;
    output n22515;
    output n73798;
    input \B_int[1] ;
    input n504;
    output n32;
    input \B_int[2] ;
    input n503;
    output \frac[26] ;
    output n30;
    input \B_int[5] ;
    input n500;
    input \addSubAB[26] ;
    input n70729;
    input \subBAExpEq[26] ;
    input n70738;
    output n33;
    input \B_int[11] ;
    input n494;
    output n37;
    input \B_int[9] ;
    input n496;
    input \B_int[14] ;
    input n491;
    input \frac[16] ;
    output n70689;
    input \B_int[17] ;
    input n488;
    output n34;
    input \B_int[16] ;
    input n489;
    output \frac[18] ;
    input \B_int[15] ;
    input n490;
    input \B_int[19] ;
    input n486;
    output n34_adj_1;
    input n70690;
    input \B_int[20] ;
    input n485;
    output n31;
    input \B_int[7] ;
    input n498;
    output \frac[10] ;
    input \B_int[21] ;
    input n484;
    input \B_int[6] ;
    input n499;
    input \B_int[3] ;
    input n502;
    output n70677;
    input \B_int[22] ;
    input n483;
    input n253;
    input n261;
    input n259;
    input n258;
    input n295;
    input n294;
    output n319;
    input n293;
    output n70658;
    input n70691;
    output \frac_sub_Norm1[25] ;
    input n356;
    output n70134;
    input n70620;
    input n70618;
    
    
    wire n10;
    wire [27:0]n243;
    wire [27:0]n272;
    
    wire n70642, n49, n70664, n70666, n70665, n68561, n114, n70651, 
        n70652, n70654, n136, n138, n67099, n6, n8, n4_c;
    wire [27:0]n330;
    
    wire n70614, n70624;
    wire [27:0]n301;
    
    wire n70619, n19020, n20382, n20380, n41796, n20588, n19016, 
        n19018, n20378, n19014, n70627, n70615, n5, n70644, n66947, 
        n66604, n21805, n70678, n70657, n70675, n105, n70648, 
        n66590, n70655, n114_adj_494, n70645, n22174, n70054, n70053, 
        n121, n70661, n70051, n70049, n70048, n70047, n66941, 
        n70649, n70686, n70684, n9, n70660, n70659, n66673, n66665, 
        n70682, n8_adj_496, n70673, n67191, n70670, n70669, n15, 
        n70653, n71720, n71721, n71722, n71723, n68777;
    
    LUT4 mux_212_i6_3_lut (.A(\A_int[28] ), .B(\B_int[28] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i6_3_lut.init = 16'hcaca;
    LUT4 mux_212_i7_3_lut (.A(\A_int[29] ), .B(\B_int[29] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i7_3_lut.init = 16'hcaca;
    LUT4 mux_212_i8_3_lut (.A(\A_int[30] ), .B(\B_int[30] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i8_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(n10), .B(\efectExp[7] ), .C(\efectExp[6] ), .D(\efectExp[5] ), 
         .Z(n62960)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 mux_53_i4_3_lut (.A(\B_int[0] ), .B(n505), .C(n61), .Z(\frac[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i4_3_lut.init = 16'hcaca;
    LUT4 mux_33_i22_3_lut (.A(\frac[21] ), .B(n70699), .C(n70634), .Z(n243[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_33_i22_3_lut.init = 16'hacac;
    LUT4 mux_33_i21_3_lut (.A(n70688), .B(n70704), .C(n70634), .Z(n243[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_33_i21_3_lut.init = 16'hacac;
    LUT4 mux_33_i20_3_lut (.A(n70687), .B(\frac[3] ), .C(n70634), .Z(n243[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_33_i20_3_lut.init = 16'hacac;
    LUT4 mux_31_i24_4_lut (.A(\frac[15] ), .B(n272[19]), .C(\leadZerosBin[2] ), 
         .D(n70634), .Z(n272[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_31_i24_4_lut.init = 16'hcac0;
    LUT4 mux_33_i24_3_lut (.A(n70681), .B(n73799), .C(n70634), .Z(n243[23])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_33_i24_3_lut.init = 16'hacac;
    LUT4 mux_31_i23_4_lut (.A(n70693), .B(n272[18]), .C(\leadZerosBin[2] ), 
         .D(n70634), .Z(n272[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_31_i23_4_lut.init = 16'hcac0;
    LUT4 mux_33_i23_3_lut (.A(n70683), .B(\frac[6] ), .C(n70634), .Z(n243[22])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_33_i23_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_4_lut (.A(\frac[3] ), .B(n70704), .C(n70642), .D(n70717), 
         .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_rep_665 (.A(\frac[3] ), .B(n70704), .C(n70642), .Z(n70635)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_665.init = 16'hfefe;
    LUT4 i1_4_lut (.A(n70664), .B(n70666), .C(n70665), .D(n68561), .Z(n114)) /* synthesis lut_function=((B ((D)+!C))+!A) */ ;
    defparam i1_4_lut.init = 16'hdd5d;
    LUT4 i1_4_lut_adj_888 (.A(n70651), .B(n70652), .C(n70654), .D(n136), 
         .Z(n138)) /* synthesis lut_function=((B ((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_888.init = 16'hdd5d;
    LUT4 i55109_2_lut (.A(\leadZerosBin[2] ), .B(n73796), .Z(n67099)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i55109_2_lut.init = 16'heeee;
    LUT4 LessThan_87_i8_3_lut_3_lut (.A(n70634), .B(\efectExp[4] ), .C(n6), 
         .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;
    defparam LessThan_87_i8_3_lut_3_lut.init = 16'he8e8;
    LUT4 LessThan_87_i6_3_lut_3_lut (.A(n73796), .B(n70782), .C(\efectExp[2] ), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;
    defparam LessThan_87_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_212_i5_3_lut (.A(\A_int[27] ), .B(\B_int[27] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i5_3_lut.init = 16'hcaca;
    LUT4 LessThan_87_i4_4_lut (.A(\efectExp[0] ), .B(\efectExp[1] ), .C(\leadZerosBin[1] ), 
         .D(\leadZerosBin[0] ), .Z(n4_c)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;
    defparam LessThan_87_i4_4_lut.init = 16'h0c8e;
    LUT4 mux_212_i3_3_lut (.A(\A_int[25] ), .B(\B_int[25] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i3_3_lut.init = 16'hcaca;
    LUT4 mux_212_i2_3_lut (.A(\A_int[24] ), .B(\B_int[24] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i2_3_lut.init = 16'hcaca;
    LUT4 mux_212_i1_3_lut (.A(\A_int[23] ), .B(\B_int[23] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i1_3_lut.init = 16'hcaca;
    LUT4 mux_22_i6_3_lut (.A(n330[5]), .B(n354), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i6_3_lut.init = 16'hcaca;
    LUT4 mux_29_i5_4_lut (.A(n296), .B(\addSubAB[0] ), .C(\leadZerosBin[2] ), 
         .D(n70617), .Z(n325)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_29_i5_4_lut.init = 16'h0aca;
    LUT4 i53968_2_lut (.A(n73796), .B(\leadZerosBin[2] ), .Z(n66873)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53968_2_lut.init = 16'heeee;
    LUT4 mux_27_i6_4_lut (.A(n70614), .B(n66873), .C(\leadZerosBin[1] ), 
         .D(n4), .Z(n330[5])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_27_i6_4_lut.init = 16'h3a0a;
    LUT4 mux_22_i8_3_lut (.A(n351), .B(n352), .C(\leadZerosBin[0] ), .Z(\frac_sub_Norm1[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i8_3_lut.init = 16'hcaca;
    LUT4 mux_22_i7_3_lut (.A(n352), .B(n330[5]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i7_3_lut.init = 16'hcaca;
    LUT4 i29350_3_lut (.A(n70634), .B(n73796), .C(n66825), .Z(n323)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29350_3_lut.init = 16'h2020;
    LUT4 mux_29_i9_4_lut (.A(n70634), .B(n296), .C(\leadZerosBin[2] ), 
         .D(n41732), .Z(n321)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_29_i9_4_lut.init = 16'hcac0;
    LUT4 i29565_4_lut (.A(n73799), .B(n70624), .C(\frac[3] ), .D(\leadZerosBin[2] ), 
         .Z(n301[7])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i29565_4_lut.init = 16'h3022;
    LUT4 mux_27_i10_3_lut (.A(n301[9]), .B(n301[7]), .C(\leadZerosBin[1] ), 
         .Z(n349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i10_3_lut.init = 16'hcaca;
    LUT4 i29351_2_lut_rep_644_3_lut (.A(n70067), .B(n70634), .C(n73796), 
         .Z(n70614)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i29351_2_lut_rep_644_3_lut.init = 16'h0808;
    LUT4 LessThan_87_i7_2_lut_rep_649_4_lut (.A(\A_int[26] ), .B(\B_int[26] ), 
         .C(\diffExpAB[8] ), .D(n73796), .Z(n70619)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam LessThan_87_i7_2_lut_rep_649_4_lut.init = 16'h35ca;
    LUT4 mux_212_i4_3_lut_rep_812 (.A(\A_int[26] ), .B(\B_int[26] ), .C(\diffExpAB[8] ), 
         .Z(n70782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i4_3_lut_rep_812.init = 16'hcaca;
    LUT4 mux_27_i12_3_lut (.A(n301[11]), .B(n301[9]), .C(\leadZerosBin[1] ), 
         .Z(n347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i12_3_lut.init = 16'hcaca;
    LUT4 mux_29_i13_3_lut (.A(n19020), .B(n41732), .C(\leadZerosBin[2] ), 
         .Z(n41774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_29_i13_3_lut.init = 16'hcaca;
    LUT4 mux_27_i14_4_lut (.A(n20382), .B(n301[11]), .C(\leadZerosBin[1] ), 
         .D(n70634), .Z(n345)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_27_i14_4_lut.init = 16'hcac0;
    LUT4 mux_27_i15_3_lut (.A(n20380), .B(n41774), .C(\leadZerosBin[1] ), 
         .Z(n41796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i15_3_lut.init = 16'hcaca;
    LUT4 mux_22_i16_3_lut (.A(n20588), .B(n41796), .C(\leadZerosBin[0] ), 
         .Z(n41812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i16_3_lut.init = 16'hcaca;
    LUT4 mux_22_i15_4_lut (.A(n70634), .B(n345), .C(\leadZerosBin[0] ), 
         .D(n41796), .Z(\frac_sub_Norm1[14] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_22_i15_4_lut.init = 16'hcac0;
    LUT4 i9039_3_lut (.A(n19016), .B(n70625), .C(\leadZerosBin[2] ), .Z(n20380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9039_3_lut.init = 16'hcaca;
    LUT4 i9041_3_lut (.A(n19018), .B(n70626), .C(\leadZerosBin[2] ), .Z(n20382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9041_3_lut.init = 16'hcaca;
    LUT4 i9243_3_lut (.A(n20378), .B(n20382), .C(\leadZerosBin[1] ), .Z(n20588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9243_3_lut.init = 16'hcaca;
    LUT4 mux_27_i17_4_lut (.A(n301[16]), .B(n20380), .C(\leadZerosBin[1] ), 
         .D(n70634), .Z(n330[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_27_i17_4_lut.init = 16'hca0a;
    LUT4 mux_22_i18_3_lut (.A(n330[17]), .B(n330[16]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i18_3_lut.init = 16'hcaca;
    LUT4 mux_22_i17_4_lut (.A(n330[16]), .B(n20588), .C(\leadZerosBin[0] ), 
         .D(n70634), .Z(\frac_sub_Norm1[16] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_22_i17_4_lut.init = 16'hca0a;
    LUT4 i7720_3_lut (.A(\frac[12] ), .B(n70704), .C(n73796), .Z(n19020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7720_3_lut.init = 16'hcaca;
    LUT4 mux_29_i17_4_lut (.A(n272[16]), .B(n19020), .C(\leadZerosBin[2] ), 
         .D(n70634), .Z(n301[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_29_i17_4_lut.init = 16'hca0a;
    LUT4 i9037_3_lut (.A(n19014), .B(n70627), .C(\leadZerosBin[2] ), .Z(n20378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9037_3_lut.init = 16'hcaca;
    LUT4 mux_27_i18_4_lut (.A(n301[17]), .B(n20378), .C(\leadZerosBin[1] ), 
         .D(n70634), .Z(n330[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_27_i18_4_lut.init = 16'hca0a;
    LUT4 mux_27_i19_3_lut (.A(n301[18]), .B(n301[16]), .C(\leadZerosBin[1] ), 
         .Z(n330[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i19_3_lut.init = 16'hcaca;
    LUT4 mux_22_i20_3_lut (.A(n330[19]), .B(n330[18]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[19] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i20_3_lut.init = 16'hcaca;
    LUT4 mux_22_i19_3_lut (.A(n330[18]), .B(n330[17]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[18] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i19_3_lut.init = 16'hcaca;
    LUT4 mux_22_i5_3_lut_4_lut (.A(n70615), .B(n70624), .C(\leadZerosBin[0] ), 
         .D(n354), .Z(\frac_sub_Norm1[4] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_22_i5_3_lut_4_lut.init = 16'h2f20;
    LUT4 i7716_3_lut (.A(n70693), .B(\frac[6] ), .C(n73796), .Z(n19016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7716_3_lut.init = 16'hcaca;
    LUT4 mux_29_i19_4_lut (.A(n272[18]), .B(n19016), .C(\leadZerosBin[2] ), 
         .D(n70634), .Z(n301[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_29_i19_4_lut.init = 16'hca0a;
    LUT4 i7718_3_lut (.A(n70692), .B(n70699), .C(n73796), .Z(n19018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7718_3_lut.init = 16'hcaca;
    LUT4 mux_29_i18_4_lut (.A(n272[17]), .B(n19018), .C(\leadZerosBin[2] ), 
         .D(n70634), .Z(n301[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_29_i18_4_lut.init = 16'hca0a;
    LUT4 mux_27_i20_3_lut (.A(n301[19]), .B(n301[17]), .C(\leadZerosBin[1] ), 
         .Z(n330[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i20_3_lut.init = 16'hcaca;
    LUT4 mux_27_i21_3_lut (.A(n301[20]), .B(n301[18]), .C(\leadZerosBin[1] ), 
         .Z(n330[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i21_3_lut.init = 16'hcaca;
    LUT4 mux_22_i22_3_lut (.A(n330[21]), .B(n330[20]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i22_3_lut.init = 16'hcaca;
    LUT4 mux_22_i21_3_lut (.A(n330[20]), .B(n330[19]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[20] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i21_3_lut.init = 16'hcaca;
    LUT4 mux_31_i17_4_lut (.A(n255), .B(n70698), .C(n73796), .D(n70634), 
         .Z(n272[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_31_i17_4_lut.init = 16'hca0a;
    LUT4 mux_29_i21_3_lut (.A(n272[20]), .B(n272[16]), .C(\leadZerosBin[2] ), 
         .Z(n301[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_29_i21_3_lut.init = 16'hcaca;
    LUT4 i7714_3_lut (.A(\frac[15] ), .B(n73799), .C(n73796), .Z(n19014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7714_3_lut.init = 16'hcaca;
    LUT4 mux_29_i20_4_lut (.A(n272[19]), .B(n19014), .C(\leadZerosBin[2] ), 
         .D(n70634), .Z(n301[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_29_i20_4_lut.init = 16'hca0a;
    LUT4 mux_27_i22_3_lut (.A(n301[21]), .B(n301[19]), .C(\leadZerosBin[1] ), 
         .Z(n330[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i22_3_lut.init = 16'hcaca;
    LUT4 mux_27_i23_3_lut (.A(n301[22]), .B(n301[20]), .C(\leadZerosBin[1] ), 
         .Z(n330[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i23_3_lut.init = 16'hcaca;
    LUT4 mux_22_i24_3_lut (.A(n330[23]), .B(n330[22]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i24_3_lut.init = 16'hcaca;
    LUT4 mux_22_i23_3_lut (.A(n330[22]), .B(n330[21]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[22] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i23_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_889 (.A(n5), .B(n70644), .C(n66947), .D(n66604), 
         .Z(n21805)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_889.init = 16'h3b33;
    LUT4 i1_4_lut_adj_890 (.A(n70635), .B(n21805), .C(n70639), .D(n73797), 
         .Z(\leadZerosBin[2] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))) */ ;
    defparam i1_4_lut_adj_890.init = 16'h8a0a;
    LUT4 mux_31_i18_4_lut (.A(n254), .B(\frac[9] ), .C(n73796), .D(n70634), 
         .Z(n272[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_31_i18_4_lut.init = 16'hca0a;
    LUT4 n10742_bdd_4_lut (.A(\leadZerosBin[2] ), .B(n70699), .C(\addSubAB[1] ), 
         .D(n70721), .Z(n70067)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam n10742_bdd_4_lut.init = 16'he444;
    LUT4 i1_4_lut_adj_891 (.A(n70678), .B(n70657), .C(n70665), .D(n70675), 
         .Z(n105)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A (B))) */ ;
    defparam i1_4_lut_adj_891.init = 16'h33b3;
    LUT4 i1_4_lut_adj_892 (.A(n105), .B(n70648), .C(n5), .D(n66604), 
         .Z(n66590)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;
    defparam i1_4_lut_adj_892.init = 16'h8c0c;
    LUT4 i1_4_lut_adj_893 (.A(n66590), .B(n70655), .C(n73797), .D(n70647), 
         .Z(n114_adj_494)) /* synthesis lut_function=(A ((C)+!B)+!A !(B ((D)+!C))) */ ;
    defparam i1_4_lut_adj_893.init = 16'hb3f3;
    LUT4 i1_4_lut_adj_894 (.A(n114_adj_494), .B(n70635), .C(n70642), .D(n70645), 
         .Z(n22174)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;
    defparam i1_4_lut_adj_894.init = 16'h8c0c;
    LUT4 i2_4_lut (.A(n22174), .B(n53), .C(n70718), .D(n49), .Z(\leadZerosBin[1] )) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i2_4_lut.init = 16'hbbbf;
    LUT4 mux_29_i22_3_lut (.A(n272[21]), .B(n272[17]), .C(\leadZerosBin[2] ), 
         .Z(n301[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_29_i22_3_lut.init = 16'hcaca;
    LUT4 i27_4_lut (.A(n70721), .B(n70054), .C(n70635), .D(n66493), 
         .Z(\leadZerosBin[0] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam i27_4_lut.init = 16'hcfc5;
    LUT4 mux_27_i24_3_lut (.A(n301[23]), .B(n301[21]), .C(\leadZerosBin[1] ), 
         .Z(n330[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_27_i24_3_lut.init = 16'hcaca;
    LUT4 mux_22_i25_3_lut (.A(n330[24]), .B(n330[23]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_22_i25_3_lut.init = 16'hcaca;
    PFUMX i55830 (.BLUT(n70053), .ALUT(n121), .C0(n70661), .Z(n70054));
    LUT4 frac_5__bdd_4_lut (.A(n70699), .B(\frac[6] ), .C(n70704), .D(n73799), 
         .Z(n70051)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam frac_5__bdd_4_lut.init = 16'hff23;
    LUT4 n70049_bdd_3_lut (.A(n70049), .B(n301[22]), .C(\leadZerosBin[1] ), 
         .Z(n330[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70049_bdd_3_lut.init = 16'hcaca;
    LUT4 n70048_bdd_3_lut (.A(n70048), .B(n272[20]), .C(\leadZerosBin[2] ), 
         .Z(n70049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70048_bdd_3_lut.init = 16'hcaca;
    PFUMX i55828 (.BLUT(n70047), .ALUT(n255), .C0(n73796), .Z(n70048));
    LUT4 n255_bdd_3_lut_56418 (.A(n70634), .B(n70680), .C(n70698), .Z(n70047)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n255_bdd_3_lut_56418.init = 16'hd8d8;
    LUT4 i1_2_lut_rep_654_4_lut_4_lut (.A(n70639), .B(n70635), .C(n66941), 
         .D(n73797), .Z(n70624)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i1_2_lut_rep_654_4_lut_4_lut.init = 16'h7fff;
    LUT4 i1_4_lut_rep_900 (.A(n70639), .B(n70635), .C(n66941), .D(n73797), 
         .Z(n73796)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;
    defparam i1_4_lut_rep_900.init = 16'h3b33;
    LUT4 i1_2_lut_rep_669_1_lut_2_lut_4_lut (.A(\B_int[4] ), .B(n501), .C(n61), 
         .D(n70649), .Z(n70639)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_669_1_lut_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_53_i8_3_lut_rep_903 (.A(\B_int[4] ), .B(n501), .C(n61), .Z(n73799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i8_3_lut_rep_903.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_1_lut_2_lut_rep_901_4_lut (.A(\B_int[8] ), .B(n497), 
         .C(n61), .D(n22515), .Z(n73797)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_3_lut_1_lut_2_lut_rep_901_4_lut.init = 16'hffca;
    LUT4 mux_53_i12_3_lut_rep_902 (.A(\B_int[8] ), .B(n497), .C(n61), 
         .Z(n73798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i12_3_lut_rep_902.init = 16'hcaca;
    LUT4 i6_2_lut_4_lut (.A(\B_int[1] ), .B(n504), .C(n61), .D(n70718), 
         .Z(n32)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i6_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_53_i5_3_lut_rep_734 (.A(\B_int[1] ), .B(n504), .C(n61), .Z(n70704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i5_3_lut_rep_734.init = 16'hcaca;
    LUT4 i5_2_lut_4_lut (.A(\B_int[2] ), .B(n503), .C(n61), .D(\frac[26] ), 
         .Z(n30)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i5_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_53_i6_3_lut_rep_729 (.A(\B_int[2] ), .B(n503), .C(n61), .Z(n70699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i6_3_lut_rep_729.init = 16'hcaca;
    LUT4 mux_53_i9_3_lut_rep_728 (.A(\B_int[5] ), .B(n500), .C(n61), .Z(n70698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i9_3_lut_rep_728.init = 16'hcaca;
    LUT4 i29457_4_lut (.A(\addSubAB[26] ), .B(n70729), .C(\subBAExpEq[26] ), 
         .D(n70738), .Z(\frac[26] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam i29457_4_lut.init = 16'heefc;
    LUT4 n70052_bdd_2_lut_3_lut (.A(n70051), .B(n70698), .C(\frac[9] ), 
         .Z(n70053)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam n70052_bdd_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i8_2_lut_4_lut (.A(\B_int[8] ), .B(n497), .C(n61), .D(n70704), 
         .Z(n33)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i8_2_lut_4_lut.init = 16'hca00;
    LUT4 i12_2_lut_4_lut (.A(\B_int[11] ), .B(n494), .C(n61), .D(\frac[9] ), 
         .Z(n37)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i12_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_53_i15_3_lut_rep_723 (.A(\B_int[11] ), .B(n494), .C(n61), 
         .Z(n70693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i15_3_lut_rep_723.init = 16'hcaca;
    LUT4 mux_53_i13_3_lut (.A(\B_int[9] ), .B(n496), .C(n61), .Z(\frac[12] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i13_3_lut.init = 16'hcaca;
    LUT4 equal_40_i17_2_lut_rep_716_4_lut (.A(\B_int[14] ), .B(n491), .C(n61), 
         .D(\frac[16] ), .Z(n70686)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam equal_40_i17_2_lut_rep_716_4_lut.init = 16'hffca;
    LUT4 mux_53_i18_3_lut_rep_719 (.A(\B_int[14] ), .B(n491), .C(n61), 
         .Z(n70689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i18_3_lut_rep_719.init = 16'hcaca;
    LUT4 i9_2_lut_4_lut (.A(\B_int[17] ), .B(n488), .C(n61), .D(\frac[15] ), 
         .Z(n34)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i9_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_53_i21_3_lut_rep_718 (.A(\B_int[17] ), .B(n488), .C(n61), 
         .Z(n70688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i21_3_lut_rep_718.init = 16'hcaca;
    LUT4 equal_55_i10_2_lut_rep_714_4_lut (.A(\B_int[16] ), .B(n489), .C(n61), 
         .D(\frac[18] ), .Z(n70684)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam equal_55_i10_2_lut_rep_714_4_lut.init = 16'hffca;
    LUT4 equal_58_i9_2_lut_4_lut (.A(\B_int[16] ), .B(n489), .C(n61), 
         .D(n70688), .Z(n9)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam equal_58_i9_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_53_i20_3_lut_rep_717 (.A(\B_int[16] ), .B(n489), .C(n61), 
         .Z(n70687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i20_3_lut_rep_717.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(\frac[16] ), .B(n70689), .C(n70660), 
         .D(n70659), .Z(n5)) /* synthesis lut_function=(A (B+(D))+!A (B+(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfecc;
    LUT4 i1_2_lut_3_lut (.A(\frac[16] ), .B(n70689), .C(\frac[15] ), .Z(n66673)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_895 (.A(\frac[18] ), .B(n70687), .C(n70688), 
         .Z(n66665)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut_adj_895.init = 16'hfefe;
    LUT4 mux_53_i19_3_lut (.A(\B_int[15] ), .B(n490), .C(n61), .Z(\frac[18] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i19_3_lut.init = 16'hcaca;
    LUT4 i8_2_lut_4_lut_adj_896 (.A(\B_int[19] ), .B(n486), .C(n61), .D(\frac[16] ), 
         .Z(n34_adj_1)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i8_2_lut_4_lut_adj_896.init = 16'hffca;
    LUT4 i1_2_lut_rep_712_4_lut (.A(\B_int[19] ), .B(n486), .C(n61), .D(\frac[21] ), 
         .Z(n70682)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_712_4_lut.init = 16'hffca;
    LUT4 mux_53_i23_3_lut_rep_713 (.A(\B_int[19] ), .B(n486), .C(n61), 
         .Z(n70683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i23_3_lut_rep_713.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut (.A(\frac[21] ), .B(n70683), .C(n66665), .Z(n8_adj_496)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'hfefe;
    LUT4 i5_4_lut (.A(n66673), .B(n70673), .C(n70690), .D(n8_adj_496), 
         .Z(n22515)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut_4_lut_adj_897 (.A(\B_int[20] ), .B(n485), .C(n61), .D(\frac[18] ), 
         .Z(n31)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i5_2_lut_4_lut_adj_897.init = 16'hffca;
    LUT4 mux_53_i11_3_lut (.A(\B_int[7] ), .B(n498), .C(n61), .Z(\frac[10] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i11_3_lut.init = 16'hcaca;
    LUT4 mux_53_i24_3_lut_rep_711 (.A(\B_int[20] ), .B(n485), .C(n61), 
         .Z(n70681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i24_3_lut_rep_711.init = 16'hcaca;
    LUT4 i1_2_lut_rep_708_4_lut (.A(\B_int[21] ), .B(n484), .C(n61), .D(n70681), 
         .Z(n70678)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_708_4_lut.init = 16'hffca;
    LUT4 mux_53_i10_3_lut (.A(\B_int[6] ), .B(n499), .C(n61), .Z(\frac[9] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i10_3_lut.init = 16'hcaca;
    LUT4 mux_53_i25_3_lut_rep_710 (.A(\B_int[21] ), .B(n484), .C(n61), 
         .Z(n70680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i25_3_lut_rep_710.init = 16'hcaca;
    LUT4 mux_53_i7_3_lut (.A(\B_int[3] ), .B(n502), .C(n61), .Z(\frac[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i7_3_lut.init = 16'hcaca;
    PFUMX LessThan_87_i10 (.BLUT(n4_c), .ALUT(n8), .C0(n67191), .Z(n10));
    LUT4 i1_2_lut_rep_703_3_lut_4_lut (.A(n70681), .B(n70680), .C(\frac[26] ), 
         .D(n70677), .Z(n70673)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_703_3_lut_4_lut.init = 16'hfffe;
    LUT4 i28185_2_lut_4_lut_3_lut (.A(n73798), .B(n22515), .C(n70639), 
         .D(n70635), .Z(n243[11])) /* synthesis lut_function=(A (C (D))) */ ;
    defparam i28185_2_lut_4_lut_3_lut.init = 16'ha000;
    LUT4 equal_76_i3_2_lut_rep_705_4_lut (.A(\B_int[22] ), .B(n483), .C(n61), 
         .D(\frac[26] ), .Z(n70675)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam equal_76_i3_2_lut_rep_705_4_lut.init = 16'hffca;
    LUT4 mux_53_i26_3_lut_rep_707 (.A(\B_int[22] ), .B(n483), .C(n61), 
         .Z(n70677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i26_3_lut_rep_707.init = 16'hcaca;
    PFUMX mux_29_i23 (.BLUT(n243[22]), .ALUT(n272[22]), .C0(n67099), .Z(n301[22]));
    PFUMX mux_29_i24 (.BLUT(n243[23]), .ALUT(n272[23]), .C0(n67099), .Z(n301[23]));
    LUT4 i1_2_lut_rep_700_3_lut_4_lut (.A(n70677), .B(\frac[26] ), .C(n70681), 
         .D(n70680), .Z(n70670)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_700_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_31_i19 (.BLUT(n253), .ALUT(n261), .C0(n73796), .Z(n272[18]));
    PFUMX mux_31_i20 (.BLUT(n243[19]), .ALUT(n243[11]), .C0(n73796), .Z(n272[19]));
    PFUMX mux_31_i21 (.BLUT(n243[20]), .ALUT(n259), .C0(n73796), .Z(n272[20]));
    PFUMX mux_31_i22 (.BLUT(n243[21]), .ALUT(n258), .C0(n73796), .Z(n272[21]));
    LUT4 i1_2_lut_rep_699_3_lut_4_lut (.A(n70677), .B(\frac[26] ), .C(n70682), 
         .D(n70678), .Z(n70669)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_699_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_29_i10 (.BLUT(n272[9]), .ALUT(n295), .C0(\leadZerosBin[2] ), 
          .Z(n301[9]));
    PFUMX mux_29_i11 (.BLUT(n272[10]), .ALUT(n294), .C0(\leadZerosBin[2] ), 
          .Z(n319));
    PFUMX mux_29_i12 (.BLUT(n272[11]), .ALUT(n293), .C0(\leadZerosBin[2] ), 
          .Z(n301[11]));
    LUT4 i1_2_lut_rep_694_3_lut_4_lut (.A(n70678), .B(n70675), .C(n70688), 
         .D(n70682), .Z(n70664)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_694_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n70678), .B(n70675), .C(n9), .D(n70682), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_696_3_lut_4_lut (.A(n70680), .B(n70675), .C(n70682), 
         .D(n70681), .Z(n70666)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_696_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_695_3_lut_4_lut (.A(n70680), .B(n70675), .C(n70683), 
         .D(n70681), .Z(n70665)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_695_3_lut_4_lut.init = 16'hfffe;
    LUT4 frac_24__bdd_4_lut (.A(n70680), .B(\frac[26] ), .C(n70681), .D(n70677), 
         .Z(n68561)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C+(D))))) */ ;
    defparam frac_24__bdd_4_lut.init = 16'h3310;
    LUT4 i28195_2_lut_rep_687_3_lut_4_lut_4_lut (.A(n70682), .B(n70673), 
         .C(n70688), .D(n70670), .Z(n70657)) /* synthesis lut_function=(A+(B (D)+!B (C (D)))) */ ;
    defparam i28195_2_lut_rep_687_3_lut_4_lut_4_lut.init = 16'hfeaa;
    LUT4 i1_2_lut_rep_691_3_lut (.A(n73798), .B(n22515), .C(\frac[10] ), 
         .Z(n70661)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_691_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_4_lut (.A(n73798), .B(n22515), .C(n138), .D(n70653), 
         .Z(n121)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B (C (D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'he222;
    LUT4 i1_2_lut_rep_685_3_lut_4_lut (.A(n73798), .B(n22515), .C(\frac[9] ), 
         .D(\frac[10] ), .Z(n70655)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_685_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_690_4_lut (.A(n70682), .B(n70670), .C(n9), .D(\frac[18] ), 
         .Z(n70660)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_690_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_689_4_lut (.A(n70683), .B(n70670), .C(\frac[21] ), 
         .D(n66665), .Z(n70659)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_689_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_688_4_lut (.A(n70688), .B(n70669), .C(n70684), .D(n66673), 
         .Z(n70658)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_688_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_679_3_lut_4_lut (.A(\frac[10] ), .B(n73797), .C(n70698), 
         .D(\frac[9] ), .Z(n70649)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_679_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_684_4_lut (.A(n70666), .B(\frac[18] ), .C(n9), .D(n70686), 
         .Z(n70654)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_684_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_682_4_lut (.A(n70666), .B(\frac[18] ), .C(n9), .D(n66673), 
         .Z(n70652)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_682_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_898 (.A(n66665), .B(\frac[21] ), .C(n70665), 
         .D(n15), .Z(n66604)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_898.init = 16'hfe00;
    LUT4 i1_2_lut_rep_683_4_lut (.A(n66673), .B(n70684), .C(n70664), .D(n70691), 
         .Z(n70653)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_683_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_681_4_lut (.A(n66673), .B(n70684), .C(n70664), .D(n70693), 
         .Z(n70651)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_681_4_lut.init = 16'hfffe;
    LUT4 i54039_3_lut_4_lut (.A(n70664), .B(n70666), .C(n70673), .D(n70665), 
         .Z(n66947)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i54039_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_675_3_lut_4_lut (.A(\frac[9] ), .B(n70661), .C(n73799), 
         .D(n70698), .Z(n70645)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_675_3_lut_4_lut.init = 16'hfffe;
    LUT4 n254_bdd_3_lut_56473 (.A(n70634), .B(n70677), .C(\frac[9] ), 
         .Z(n71720)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n254_bdd_3_lut_56473.init = 16'hd8d8;
    LUT4 i1_4_lut_4_lut_adj_899 (.A(n70689), .B(n70659), .C(n114), .D(n15), 
         .Z(n136)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B (C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_899.init = 16'he222;
    PFUMX i56469 (.BLUT(n71720), .ALUT(n254), .C0(n73796), .Z(n71721));
    LUT4 n71721_bdd_3_lut (.A(n71721), .B(n272[21]), .C(\leadZerosBin[2] ), 
         .Z(n71722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n71721_bdd_3_lut.init = 16'hcaca;
    LUT4 n71722_bdd_3_lut (.A(n71722), .B(n301[23]), .C(\leadZerosBin[1] ), 
         .Z(n71723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n71722_bdd_3_lut.init = 16'hcaca;
    PFUMX i56471 (.BLUT(n71723), .ALUT(n330[24]), .C0(\leadZerosBin[0] ), 
          .Z(\frac_sub_Norm1[25] ));
    LUT4 i1_2_lut_rep_678_3_lut_4_lut (.A(n66673), .B(n70660), .C(n70658), 
         .D(n70693), .Z(n70648)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_678_3_lut_4_lut.init = 16'heee0;
    LUT4 i1_2_lut_rep_674_3_lut_4_lut (.A(n70652), .B(n70651), .C(n22515), 
         .D(n70653), .Z(n70644)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_674_3_lut_4_lut.init = 16'h8000;
    LUT4 i29358_2_lut_4_lut (.A(n73798), .B(\frac[3] ), .C(n73796), .D(n70634), 
         .Z(n272[11])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29358_2_lut_4_lut.init = 16'hca00;
    LUT4 i1_3_lut_rep_672_4_lut (.A(n73799), .B(n70649), .C(\frac[6] ), 
         .D(n70699), .Z(n70642)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_rep_672_4_lut.init = 16'hfffe;
    LUT4 i7722_3_lut_rep_657 (.A(n73798), .B(\frac[3] ), .C(n73796), .Z(n70627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7722_3_lut_rep_657.init = 16'hcaca;
    LUT4 i54033_3_lut_4_lut (.A(n70647), .B(n70648), .C(n5), .D(n66604), 
         .Z(n66941)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i54033_3_lut_4_lut.init = 16'h8000;
    LUT4 leadZerosBin_1__bdd_4_lut_56072 (.A(\leadZerosBin[1] ), .B(\frac[3] ), 
         .C(\addSubAB[1] ), .D(n70721), .Z(n68777)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam leadZerosBin_1__bdd_4_lut_56072.init = 16'he444;
    LUT4 n6_bdd_3_lut_4_lut (.A(n70615), .B(n70624), .C(\leadZerosBin[0] ), 
         .D(n356), .Z(n70134)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;
    defparam n6_bdd_3_lut_4_lut.init = 16'hf202;
    LUT4 i2_3_lut_rep_664_4_lut (.A(n70645), .B(n70642), .C(n70635), .D(n73797), 
         .Z(n70634)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_664_4_lut.init = 16'h8000;
    LUT4 i29360_2_lut_4_lut (.A(\frac[9] ), .B(n70718), .C(n73796), .D(n70634), 
         .Z(n272[9])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29360_2_lut_4_lut.init = 16'hca00;
    LUT4 i29359_2_lut_4_lut (.A(\frac[10] ), .B(n70717), .C(n73796), .D(n70634), 
         .Z(n272[10])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29359_2_lut_4_lut.init = 16'hca00;
    LUT4 i55077_4_lut_4_lut (.A(n70620), .B(\efectExp[2] ), .C(\leadZerosBin[2] ), 
         .D(n70619), .Z(n67191)) /* synthesis lut_function=((B ((D)+!C)+!B (C+(D)))+!A) */ ;
    defparam i55077_4_lut_4_lut.init = 16'hff7d;
    LUT4 n68777_bdd_2_lut_rep_645 (.A(n68777), .B(\leadZerosBin[2] ), .Z(n70615)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n68777_bdd_2_lut_rep_645.init = 16'h2222;
    LUT4 mux_27_i8_3_lut_4_lut (.A(n70618), .B(n73796), .C(\leadZerosBin[1] ), 
         .D(n301[7]), .Z(n351)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_27_i8_3_lut_4_lut.init = 16'h2f20;
    
endmodule
//
// Verilog Description of module \right_shifter(27,8,4) 
//

module \right_shifter(27,8,4)  (diffExpAB, diffExpBA, \diffExp[4] , n70763, 
            \B_int[21] , \A_int[21] , \diffExp[1] , \B_int[19] , \A_int[19] , 
            \B_int[14] , \A_int[14] , \B_int[15] , \A_int[15] , \B_int[13] , 
            \A_int[13] , \B_int[7] , \A_int[7] , \B_int[4] , \A_int[4] , 
            \efectFracB[13] , \diffExp[2] , n70734, n15, \efectFracB[15] , 
            \efectFracB[14] , \fracAlign_int[0] , n7, \efectFracB_align[2] , 
            \efectFracB_align[1] , \B_int[0] , \A_int[0] , \B_int[1] , 
            \A_int[1] , \fracAlign_int[4] , \fracAlign_int[3] , \B_int[3] , 
            \A_int[3] , \B_int[2] , \A_int[2] , \fracAlign_int[6] , 
            \fracAlign_int[5] , \B_int[5] , \A_int[5] , \fracAlign_int[8] , 
            \fracAlign_int[7] , \B_int[6] , \A_int[6] , \fracAlign_int[10] , 
            \fracAlign_int[9] , \B_int[9] , \A_int[9] , \B_int[8] , 
            \A_int[8] , \fracAlign_int[12] , n66898, n41776, \fracAlign_int[14] , 
            \fracAlign_int[13] , \fracAlign_int[16] , \fracAlign_int[15] , 
            \fracAlign_int[18] , \fracAlign_int[17] , \B_int[17] , \A_int[17] , 
            \B_int[16] , \A_int[16] , \B_int[18] , \A_int[18] , \fracAlign_int[20] , 
            n41584, \fracAlign_int[22] , \fracAlign_int[21] , \B_int[20] , 
            \A_int[20] , n66912, \B_int[22] , \A_int[22] , n66221, 
            n458, n70727, n61, \frac[21] , n463, \frac[16] );
    input [8:0]diffExpAB;
    input [8:0]diffExpBA;
    output \diffExp[4] ;
    output n70763;
    input \B_int[21] ;
    input \A_int[21] ;
    output \diffExp[1] ;
    input \B_int[19] ;
    input \A_int[19] ;
    input \B_int[14] ;
    input \A_int[14] ;
    input \B_int[15] ;
    input \A_int[15] ;
    input \B_int[13] ;
    input \A_int[13] ;
    input \B_int[7] ;
    input \A_int[7] ;
    input \B_int[4] ;
    input \A_int[4] ;
    input \efectFracB[13] ;
    output \diffExp[2] ;
    output n70734;
    output n15;
    input \efectFracB[15] ;
    input \efectFracB[14] ;
    output \fracAlign_int[0] ;
    output n7;
    output \efectFracB_align[2] ;
    output \efectFracB_align[1] ;
    input \B_int[0] ;
    input \A_int[0] ;
    input \B_int[1] ;
    input \A_int[1] ;
    output \fracAlign_int[4] ;
    output \fracAlign_int[3] ;
    input \B_int[3] ;
    input \A_int[3] ;
    input \B_int[2] ;
    input \A_int[2] ;
    output \fracAlign_int[6] ;
    output \fracAlign_int[5] ;
    input \B_int[5] ;
    input \A_int[5] ;
    output \fracAlign_int[8] ;
    output \fracAlign_int[7] ;
    input \B_int[6] ;
    input \A_int[6] ;
    output \fracAlign_int[10] ;
    output \fracAlign_int[9] ;
    input \B_int[9] ;
    input \A_int[9] ;
    input \B_int[8] ;
    input \A_int[8] ;
    output \fracAlign_int[12] ;
    output n66898;
    output n41776;
    output \fracAlign_int[14] ;
    output \fracAlign_int[13] ;
    output \fracAlign_int[16] ;
    output \fracAlign_int[15] ;
    output \fracAlign_int[18] ;
    output \fracAlign_int[17] ;
    input \B_int[17] ;
    input \A_int[17] ;
    input \B_int[16] ;
    input \A_int[16] ;
    input \B_int[18] ;
    input \A_int[18] ;
    output \fracAlign_int[20] ;
    output n41584;
    output \fracAlign_int[22] ;
    output \fracAlign_int[21] ;
    input \B_int[20] ;
    input \A_int[20] ;
    output n66912;
    input \B_int[22] ;
    input \A_int[22] ;
    output n66221;
    input n458;
    input n70727;
    input n61;
    output \frac[21] ;
    input n463;
    output \frac[16] ;
    
    wire [27:0]efectFracB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(67[23:33])
    wire [8:0]diffExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[33:40])
    
    wire n70803, n70762, n70802, n70801, n70756, n70800, n70755, 
        n70799, n70747, n70798, n70757, n70797, n16, n70796;
    wire [27:0]n37;
    
    wire n28, n66597;
    wire [27:0]n69;
    
    wire n70761, n20394, n41432, n19106, n41654, n70760, n70759, 
        n70758, n70732;
    wire [27:0]n5;
    
    wire n14, n13, n6, n19820, n66881, n66883, n22, n20, n24_adj_491, 
        n17503;
    wire [27:0]n101;
    
    wire n67021, n63125, n19110, n19112, n19108, n20402, n20400, 
        n20596, n20398, n41734, n20396, n20594, n23577, n35487, 
        n35482, n70872, n70873;
    
    LUT4 i28984_2_lut_rep_793_4_lut (.A(diffExpAB[3]), .B(diffExpBA[3]), 
         .C(diffExpAB[8]), .D(\diffExp[4] ), .Z(n70763)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i28984_2_lut_rep_793_4_lut.init = 16'hffca;
    LUT4 mux_2994_i4_3_lut_rep_833 (.A(diffExpAB[3]), .B(diffExpBA[3]), 
         .C(diffExpAB[8]), .Z(n70803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2994_i4_3_lut_rep_833.init = 16'hcaca;
    LUT4 i1_2_lut_rep_792_4_lut (.A(\B_int[21] ), .B(\A_int[21] ), .C(diffExpAB[8]), 
         .D(\diffExp[1] ), .Z(n70762)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_792_4_lut.init = 16'hffca;
    LUT4 mux_3878_i22_3_lut_rep_832 (.A(\B_int[21] ), .B(\A_int[21] ), .C(diffExpAB[8]), 
         .Z(n70802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i22_3_lut_rep_832.init = 16'hcaca;
    LUT4 mux_3878_i20_3_lut_rep_831 (.A(\B_int[19] ), .B(\A_int[19] ), .C(diffExpAB[8]), 
         .Z(n70801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i20_3_lut_rep_831.init = 16'hcaca;
    LUT4 i1_2_lut_rep_786_4_lut (.A(\B_int[14] ), .B(\A_int[14] ), .C(diffExpAB[8]), 
         .D(\diffExp[4] ), .Z(n70756)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_786_4_lut.init = 16'hca00;
    LUT4 i23870_3_lut_rep_830 (.A(\B_int[14] ), .B(\A_int[14] ), .C(diffExpAB[8]), 
         .Z(n70800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23870_3_lut_rep_830.init = 16'hcaca;
    LUT4 i28238_2_lut_rep_785_4_lut (.A(\B_int[15] ), .B(\A_int[15] ), .C(diffExpAB[8]), 
         .D(\diffExp[4] ), .Z(n70755)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i28238_2_lut_rep_785_4_lut.init = 16'hca00;
    LUT4 mux_3878_i16_3_lut_rep_829 (.A(\B_int[15] ), .B(\A_int[15] ), .C(diffExpAB[8]), 
         .Z(n70799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i16_3_lut_rep_829.init = 16'hcaca;
    LUT4 i1_2_lut_rep_777_4_lut (.A(\B_int[13] ), .B(\A_int[13] ), .C(diffExpAB[8]), 
         .D(\diffExp[4] ), .Z(n70747)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_777_4_lut.init = 16'hca00;
    LUT4 i23883_3_lut_rep_828 (.A(\B_int[13] ), .B(\A_int[13] ), .C(diffExpAB[8]), 
         .Z(n70798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23883_3_lut_rep_828.init = 16'hcaca;
    LUT4 i28237_2_lut_rep_787_4_lut (.A(\B_int[7] ), .B(\A_int[7] ), .C(diffExpAB[8]), 
         .D(\diffExp[4] ), .Z(n70757)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i28237_2_lut_rep_787_4_lut.init = 16'hffca;
    LUT4 mux_3878_i8_3_lut_rep_827 (.A(\B_int[7] ), .B(\A_int[7] ), .C(diffExpAB[8]), 
         .Z(n70797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i8_3_lut_rep_827.init = 16'hcaca;
    LUT4 i3_2_lut_4_lut (.A(\B_int[4] ), .B(\A_int[4] ), .C(diffExpAB[8]), 
         .D(\efectFracB[13] ), .Z(n16)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i3_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_3878_i5_3_lut_rep_826 (.A(\B_int[4] ), .B(\A_int[4] ), .C(diffExpAB[8]), 
         .Z(n70796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i5_3_lut_rep_826.init = 16'hcaca;
    LUT4 i29375_2_lut_3_lut (.A(\diffExp[4] ), .B(n70803), .C(n70801), 
         .Z(n37[22])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29375_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut (.A(\diffExp[4] ), .B(n70803), .C(efectFracB[21]), 
         .Z(n28)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i29376_2_lut_3_lut (.A(\diffExp[4] ), .B(n70803), .C(efectFracB[20]), 
         .Z(n37[20])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29376_2_lut_3_lut.init = 16'h1010;
    LUT4 i29377_2_lut_3_lut (.A(\diffExp[4] ), .B(n70803), .C(efectFracB[19]), 
         .Z(n37[19])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29377_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\diffExp[4] ), .B(n70803), .C(n70801), 
         .D(\diffExp[2] ), .Z(n66597)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i29573_2_lut_3_lut_4_lut (.A(\diffExp[4] ), .B(n70803), .C(n70802), 
         .D(\diffExp[2] ), .Z(n69[24])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i29573_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i29574_2_lut_3_lut_4_lut (.A(\diffExp[4] ), .B(n70803), .C(efectFracB[23]), 
         .D(\diffExp[2] ), .Z(n69[23])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i29574_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i2_2_lut_rep_764_3_lut (.A(\diffExp[4] ), .B(n70803), .C(\diffExp[2] ), 
         .Z(n70734)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_2_lut_rep_764_3_lut.init = 16'hfefe;
    LUT4 i24_4_lut_4_lut (.A(n70802), .B(\diffExp[1] ), .C(diffExp[0]), 
         .D(efectFracB[25]), .Z(n15)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam i24_4_lut_4_lut.init = 16'h3e0e;
    LUT4 i29627_2_lut_4_lut (.A(efectFracB[21]), .B(efectFracB[25]), .C(\diffExp[2] ), 
         .D(n70763), .Z(n69[21])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29627_2_lut_4_lut.init = 16'h00ca;
    LUT4 i9051_3_lut_rep_791 (.A(efectFracB[21]), .B(efectFracB[25]), .C(\diffExp[2] ), 
         .Z(n70761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9051_3_lut_rep_791.init = 16'hcaca;
    LUT4 i9047_3_lut_4_lut (.A(\diffExp[2] ), .B(n70801), .C(\diffExp[1] ), 
         .D(n20394), .Z(n41432)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i9047_3_lut_4_lut.init = 16'hefe0;
    LUT4 i29841_2_lut_3_lut (.A(n70803), .B(n70799), .C(\diffExp[4] ), 
         .Z(n37[18])) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i29841_2_lut_3_lut.init = 16'h0e0e;
    LUT4 mux_3928_i15_3_lut_4_lut (.A(n70803), .B(n70799), .C(\diffExp[2] ), 
         .D(n19106), .Z(n41654)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3928_i15_3_lut_4_lut.init = 16'hefe0;
    LUT4 i29378_2_lut_4_lut (.A(n70800), .B(efectFracB[25]), .C(n70803), 
         .D(\diffExp[4] ), .Z(n37[17])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29378_2_lut_4_lut.init = 16'h00ca;
    LUT4 i7800_3_lut_rep_790 (.A(n70800), .B(efectFracB[25]), .C(n70803), 
         .Z(n70760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7800_3_lut_rep_790.init = 16'hcaca;
    LUT4 i29380_2_lut_4_lut (.A(\efectFracB[15] ), .B(efectFracB[23]), .C(n70803), 
         .D(\diffExp[4] ), .Z(n37[15])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29380_2_lut_4_lut.init = 16'h00ca;
    LUT4 i7804_3_lut_rep_789 (.A(\efectFracB[15] ), .B(efectFracB[23]), 
         .C(n70803), .Z(n70759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7804_3_lut_rep_789.init = 16'hcaca;
    LUT4 i29379_2_lut_4_lut (.A(n70798), .B(n70802), .C(n70803), .D(\diffExp[4] ), 
         .Z(n37[16])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29379_2_lut_4_lut.init = 16'h00ca;
    LUT4 i7802_3_lut_rep_788 (.A(n70798), .B(n70802), .C(n70803), .Z(n70758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7802_3_lut_rep_788.init = 16'hcaca;
    LUT4 mux_3923_i3_3_lut_rep_762_4_lut_4_lut (.A(n70797), .B(\diffExp[4] ), 
         .C(n70803), .D(n70799), .Z(n70732)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;
    defparam mux_3923_i3_3_lut_rep_762_4_lut_4_lut.init = 16'hece0;
    LUT4 mux_3923_i11_4_lut_4_lut (.A(n70797), .B(\diffExp[4] ), .C(n70803), 
         .D(n70799), .Z(n37[10])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam mux_3923_i11_4_lut_4_lut.init = 16'h3e0e;
    LUT4 mux_3923_i2_3_lut_4_lut (.A(\diffExp[4] ), .B(n70800), .C(n70803), 
         .D(n5[9]), .Z(n37[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_3923_i2_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_3923_i1_3_lut_4_lut (.A(\diffExp[4] ), .B(n70798), .C(n70803), 
         .D(n5[8]), .Z(n37[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_3923_i1_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_3928_i1_3_lut (.A(n37[0]), .B(n37[4]), .C(\diffExp[2] ), 
         .Z(n69[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i1_3_lut.init = 16'hcaca;
    LUT4 i6_4_lut (.A(n5[6]), .B(n5[3]), .C(n5[4]), .D(n70747), .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i5_4_lut (.A(n5[7]), .B(n70756), .C(n70755), .D(n5[5]), .Z(n13)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i8518_4_lut (.A(\diffExp[2] ), .B(n37[0]), .C(n6), .D(n37[1]), 
         .Z(n19820)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i8518_4_lut.init = 16'haaa8;
    LUT4 i53976_3_lut (.A(\diffExp[1] ), .B(n69[0]), .C(n69[1]), .Z(n66881)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i53976_3_lut.init = 16'ha8a8;
    LUT4 i53978_4_lut (.A(n69[0]), .B(n19820), .C(n69[2]), .D(\diffExp[1] ), 
         .Z(n66883)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i53978_4_lut.init = 16'hfcee;
    LUT4 i9_4_lut (.A(n70797), .B(\efectFracB[14] ), .C(efectFracB[3]), 
         .D(efectFracB[6]), .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_3_lut (.A(efectFracB[4]), .B(efectFracB[11]), .C(efectFracB[12]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i11_4_lut (.A(\efectFracB[15] ), .B(n22), .C(n16), .D(efectFracB[8]), 
         .Z(n24_adj_491)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i6859_3_lut (.A(n13), .B(n70803), .C(n14), .Z(n17503)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i6859_3_lut.init = 16'hc8c8;
    LUT4 i54110_4_lut (.A(n101[1]), .B(n66883), .C(n66881), .D(diffExp[0]), 
         .Z(n67021)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i54110_4_lut.init = 16'hfefc;
    LUT4 i12_4_lut (.A(efectFracB[5]), .B(n24_adj_491), .C(n20), .D(efectFracB[9]), 
         .Z(n63125)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i54122_4_lut (.A(n63125), .B(n67021), .C(n17503), .D(\diffExp[4] ), 
         .Z(\fracAlign_int[0] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i54122_4_lut.init = 16'hfefc;
    LUT4 mux_3928_i3_3_lut (.A(n70732), .B(n37[6]), .C(\diffExp[2] ), 
         .Z(n69[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i3_3_lut.init = 16'hcaca;
    LUT4 mux_3928_i2_3_lut (.A(n37[1]), .B(n37[5]), .C(\diffExp[2] ), 
         .Z(n69[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i2_3_lut (.A(n69[1]), .B(n69[3]), .C(\diffExp[1] ), 
         .Z(n101[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i3_3_lut (.A(n69[2]), .B(n69[4]), .C(\diffExp[1] ), 
         .Z(n101[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i3_3_lut.init = 16'hcaca;
    LUT4 i28220_4_lut (.A(n101[2]), .B(n7), .C(n101[3]), .D(diffExp[0]), 
         .Z(\efectFracB_align[2] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i28220_4_lut.init = 16'h3022;
    LUT4 i28221_4_lut (.A(n101[1]), .B(n7), .C(n101[2]), .D(diffExp[0]), 
         .Z(\efectFracB_align[1] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i28221_4_lut.init = 16'h3022;
    LUT4 mux_3878_i1_3_lut (.A(\B_int[0] ), .B(\A_int[0] ), .C(diffExpAB[8]), 
         .Z(efectFracB[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i1_3_lut.init = 16'hcaca;
    LUT4 mux_3918_i4_3_lut (.A(efectFracB[3]), .B(efectFracB[19]), .C(\diffExp[4] ), 
         .Z(n5[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3918_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i4_4_lut (.A(n5[3]), .B(efectFracB[11]), .C(n70803), 
         .D(\diffExp[4] ), .Z(n37[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3923_i4_4_lut.init = 16'h0aca;
    LUT4 mux_3928_i4_3_lut (.A(n37[3]), .B(n37[7]), .C(\diffExp[2] ), 
         .Z(n69[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i4_3_lut (.A(n69[3]), .B(n69[5]), .C(\diffExp[1] ), 
         .Z(n101[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i2_3_lut (.A(\B_int[1] ), .B(\A_int[1] ), .C(diffExpAB[8]), 
         .Z(efectFracB[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3918_i5_3_lut (.A(efectFracB[4]), .B(efectFracB[20]), .C(\diffExp[4] ), 
         .Z(n5[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3918_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i5_4_lut (.A(n5[4]), .B(efectFracB[12]), .C(n70803), 
         .D(\diffExp[4] ), .Z(n37[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3923_i5_4_lut.init = 16'h0aca;
    LUT4 mux_3928_i5_3_lut (.A(n37[4]), .B(n37[8]), .C(\diffExp[2] ), 
         .Z(n69[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i5_3_lut (.A(n69[4]), .B(n69[6]), .C(\diffExp[1] ), 
         .Z(n101[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i5_3_lut (.A(n101[4]), .B(n101[5]), .C(diffExp[0]), 
         .Z(\fracAlign_int[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i4_3_lut (.A(n101[3]), .B(n101[4]), .C(diffExp[0]), 
         .Z(\fracAlign_int[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i4_3_lut (.A(\B_int[3] ), .B(\A_int[3] ), .C(diffExpAB[8]), 
         .Z(efectFracB[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3918_i7_3_lut (.A(efectFracB[6]), .B(n70801), .C(\diffExp[4] ), 
         .Z(n5[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3918_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i7_4_lut (.A(n5[6]), .B(\diffExp[4] ), .C(n70803), .D(\efectFracB[14] ), 
         .Z(n37[6])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3923_i7_4_lut.init = 16'h3a0a;
    LUT4 mux_3928_i7_3_lut (.A(n37[6]), .B(n37[10]), .C(\diffExp[2] ), 
         .Z(n69[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i3_3_lut (.A(\B_int[2] ), .B(\A_int[2] ), .C(diffExpAB[8]), 
         .Z(efectFracB[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i3_3_lut.init = 16'hcaca;
    LUT4 i12_3_lut (.A(efectFracB[5]), .B(efectFracB[21]), .C(\diffExp[4] ), 
         .Z(n5[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i6_4_lut (.A(n5[5]), .B(\diffExp[4] ), .C(n70803), .D(\efectFracB[13] ), 
         .Z(n37[5])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3923_i6_4_lut.init = 16'h3a0a;
    LUT4 mux_3928_i6_3_lut (.A(n37[5]), .B(n37[9]), .C(\diffExp[2] ), 
         .Z(n69[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3928_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i6_3_lut (.A(n69[5]), .B(n69[7]), .C(\diffExp[1] ), 
         .Z(n101[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i7_3_lut (.A(n69[6]), .B(n69[8]), .C(\diffExp[1] ), 
         .Z(n101[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i7_3_lut (.A(n101[6]), .B(n101[7]), .C(diffExp[0]), 
         .Z(\fracAlign_int[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i6_3_lut (.A(n101[5]), .B(n101[6]), .C(diffExp[0]), 
         .Z(\fracAlign_int[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i6_3_lut (.A(\B_int[5] ), .B(\A_int[5] ), .C(diffExpAB[8]), 
         .Z(efectFracB[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3918_i9_3_lut (.A(efectFracB[8]), .B(n70802), .C(\diffExp[4] ), 
         .Z(n5[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3918_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i9_4_lut (.A(n5[8]), .B(\diffExp[4] ), .C(n70803), .D(n70798), 
         .Z(n37[8])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3923_i9_4_lut.init = 16'h3a0a;
    LUT4 mux_3928_i9_4_lut (.A(n37[8]), .B(n19110), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3928_i9_4_lut.init = 16'h0aca;
    LUT4 mux_3918_i8_3_lut (.A(n70796), .B(efectFracB[23]), .C(\diffExp[4] ), 
         .Z(n5[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3918_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i8_4_lut (.A(n5[7]), .B(\efectFracB[15] ), .C(n70803), 
         .D(\diffExp[4] ), .Z(n37[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3923_i8_4_lut.init = 16'h0aca;
    LUT4 mux_3928_i8_4_lut (.A(n37[7]), .B(n19112), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3928_i8_4_lut.init = 16'h0aca;
    LUT4 mux_3933_i8_3_lut (.A(n69[7]), .B(n69[9]), .C(\diffExp[1] ), 
         .Z(n101[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i9_3_lut (.A(n69[8]), .B(n69[10]), .C(\diffExp[1] ), 
         .Z(n101[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i9_3_lut (.A(n101[8]), .B(n101[9]), .C(diffExp[0]), 
         .Z(\fracAlign_int[8] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i8_3_lut (.A(n101[7]), .B(n101[8]), .C(diffExp[0]), 
         .Z(\fracAlign_int[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3928_i11_4_lut (.A(n37[10]), .B(n19106), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3928_i11_4_lut.init = 16'h0aca;
    LUT4 mux_3878_i7_3_lut (.A(\B_int[6] ), .B(\A_int[6] ), .C(diffExpAB[8]), 
         .Z(efectFracB[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3918_i10_3_lut (.A(efectFracB[9]), .B(efectFracB[25]), .C(\diffExp[4] ), 
         .Z(n5[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3918_i10_3_lut.init = 16'hcaca;
    LUT4 mux_3923_i10_4_lut (.A(n5[9]), .B(\diffExp[4] ), .C(n70803), 
         .D(n70800), .Z(n37[9])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3923_i10_4_lut.init = 16'h3a0a;
    LUT4 mux_3928_i10_4_lut (.A(n37[9]), .B(n19108), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3928_i10_4_lut.init = 16'h0aca;
    LUT4 mux_3933_i10_4_lut (.A(n69[9]), .B(n20402), .C(\diffExp[1] ), 
         .D(\diffExp[4] ), .Z(n101[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3933_i10_4_lut.init = 16'h0aca;
    LUT4 mux_3933_i11_4_lut (.A(n69[10]), .B(n20400), .C(\diffExp[1] ), 
         .D(\diffExp[4] ), .Z(n101[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3933_i11_4_lut.init = 16'h0aca;
    LUT4 mux_3938_i11_4_lut (.A(n101[10]), .B(n20596), .C(diffExp[0]), 
         .D(\diffExp[4] ), .Z(\fracAlign_int[10] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3938_i11_4_lut.init = 16'h0aca;
    LUT4 mux_3938_i10_3_lut (.A(n101[9]), .B(n101[10]), .C(diffExp[0]), 
         .Z(\fracAlign_int[9] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i10_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i10_3_lut (.A(\B_int[9] ), .B(\A_int[9] ), .C(diffExpAB[8]), 
         .Z(efectFracB[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i10_3_lut.init = 16'hcaca;
    LUT4 i7810_3_lut (.A(efectFracB[12]), .B(efectFracB[20]), .C(n70803), 
         .Z(n19110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7810_3_lut.init = 16'hcaca;
    LUT4 i9059_3_lut (.A(n19110), .B(n70758), .C(\diffExp[2] ), .Z(n20400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9059_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i9_3_lut (.A(\B_int[8] ), .B(\A_int[8] ), .C(diffExpAB[8]), 
         .Z(efectFracB[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i9_3_lut.init = 16'hcaca;
    LUT4 i7812_3_lut (.A(efectFracB[11]), .B(efectFracB[19]), .C(n70803), 
         .Z(n19112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7812_3_lut.init = 16'hcaca;
    LUT4 i9061_3_lut (.A(n19112), .B(n70759), .C(\diffExp[2] ), .Z(n20402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9061_3_lut.init = 16'hcaca;
    LUT4 i9251_3_lut (.A(n20402), .B(n20398), .C(\diffExp[1] ), .Z(n20596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9251_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i13_3_lut (.A(n20400), .B(n41654), .C(\diffExp[1] ), 
         .Z(n41734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i13_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i13_4_lut (.A(\diffExp[4] ), .B(n101[13]), .C(diffExp[0]), 
         .D(n41734), .Z(\fracAlign_int[12] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3938_i13_4_lut.init = 16'hc5c0;
    LUT4 i53992_3_lut_4_lut (.A(\diffExp[2] ), .B(n70763), .C(efectFracB[25]), 
         .D(diffExp[0]), .Z(n66898)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i53992_3_lut_4_lut.init = 16'h1110;
    LUT4 mux_3938_i12_3_lut (.A(n20596), .B(n41734), .C(diffExp[0]), .Z(n41776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i12_3_lut.init = 16'hcaca;
    LUT4 i7808_3_lut (.A(\efectFracB[13] ), .B(efectFracB[21]), .C(n70803), 
         .Z(n19108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7808_3_lut.init = 16'hcaca;
    LUT4 i9057_3_lut (.A(n19108), .B(n70760), .C(\diffExp[2] ), .Z(n20398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9057_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i14_4_lut (.A(n20398), .B(n69[15]), .C(\diffExp[1] ), 
         .D(\diffExp[4] ), .Z(n101[13])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam mux_3933_i14_4_lut.init = 16'hc0ca;
    LUT4 i2_2_lut_4_lut (.A(n70755), .B(n70757), .C(n70803), .D(n37[3]), 
         .Z(n6)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i2_2_lut_4_lut.init = 16'hffca;
    LUT4 i7806_3_lut (.A(\efectFracB[14] ), .B(n70801), .C(n70803), .Z(n19106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7806_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i15_4_lut (.A(\diffExp[4] ), .B(n69[16]), .C(\diffExp[1] ), 
         .D(n41654), .Z(n101[14])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3933_i15_4_lut.init = 16'hc5c0;
    LUT4 mux_3938_i15_3_lut (.A(n101[14]), .B(n101[15]), .C(diffExp[0]), 
         .Z(\fracAlign_int[14] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i15_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i14_3_lut (.A(n101[13]), .B(n101[14]), .C(diffExp[0]), 
         .Z(\fracAlign_int[13] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i14_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i16_3_lut (.A(n69[15]), .B(n69[17]), .C(\diffExp[1] ), 
         .Z(n101[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i16_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i17_3_lut (.A(n69[16]), .B(n69[18]), .C(\diffExp[1] ), 
         .Z(n101[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3933_i17_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i17_3_lut (.A(n101[16]), .B(n101[17]), .C(diffExp[0]), 
         .Z(\fracAlign_int[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i17_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i16_3_lut (.A(n101[15]), .B(n101[16]), .C(diffExp[0]), 
         .Z(\fracAlign_int[15] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i16_3_lut.init = 16'hcaca;
    LUT4 mux_3933_i18_4_lut (.A(n69[17]), .B(n20396), .C(\diffExp[1] ), 
         .D(n70763), .Z(n101[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3933_i18_4_lut.init = 16'h0aca;
    LUT4 mux_3933_i19_4_lut (.A(n69[18]), .B(n20394), .C(\diffExp[1] ), 
         .D(n70763), .Z(n101[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3933_i19_4_lut.init = 16'h0aca;
    LUT4 mux_3938_i19_4_lut (.A(n101[18]), .B(n20594), .C(diffExp[0]), 
         .D(n70763), .Z(\fracAlign_int[18] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3938_i19_4_lut.init = 16'h0aca;
    LUT4 mux_3938_i18_3_lut (.A(n101[17]), .B(n101[18]), .C(diffExp[0]), 
         .Z(\fracAlign_int[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i18_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i18_3_lut (.A(\B_int[17] ), .B(\A_int[17] ), .C(diffExpAB[8]), 
         .Z(efectFracB[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i18_3_lut.init = 16'hcaca;
    LUT4 i9053_3_lut (.A(efectFracB[20]), .B(n70802), .C(\diffExp[2] ), 
         .Z(n20394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9053_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i17_3_lut (.A(\B_int[16] ), .B(\A_int[16] ), .C(diffExpAB[8]), 
         .Z(efectFracB[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i17_3_lut.init = 16'hcaca;
    LUT4 i23865_3_lut (.A(\B_int[18] ), .B(\A_int[18] ), .C(diffExpAB[8]), 
         .Z(efectFracB[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23865_3_lut.init = 16'hcaca;
    LUT4 i9055_3_lut (.A(efectFracB[19]), .B(efectFracB[23]), .C(\diffExp[2] ), 
         .Z(n20396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9055_3_lut.init = 16'hcaca;
    LUT4 i9249_3_lut (.A(n20396), .B(n70761), .C(\diffExp[1] ), .Z(n20594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9249_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i21_4_lut (.A(n41432), .B(n101[21]), .C(diffExp[0]), 
         .D(n70763), .Z(\fracAlign_int[20] )) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam mux_3938_i21_4_lut.init = 16'hc0ca;
    LUT4 i9247_3_lut (.A(n20594), .B(n41432), .C(diffExp[0]), .Z(n41584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9247_3_lut.init = 16'hcaca;
    LUT4 mux_3938_i23_4_lut (.A(n101[22]), .B(n23577), .C(diffExp[0]), 
         .D(n70734), .Z(\fracAlign_int[22] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3938_i23_4_lut.init = 16'h0aca;
    LUT4 mux_3938_i22_3_lut (.A(n101[21]), .B(n101[22]), .C(diffExp[0]), 
         .Z(\fracAlign_int[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3938_i22_3_lut.init = 16'hcaca;
    LUT4 mux_3878_i21_3_lut (.A(\B_int[20] ), .B(\A_int[20] ), .C(diffExpAB[8]), 
         .Z(efectFracB[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i21_3_lut.init = 16'hcaca;
    LUT4 i11894_3_lut (.A(efectFracB[23]), .B(efectFracB[25]), .C(\diffExp[1] ), 
         .Z(n23577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11894_3_lut.init = 16'hcaca;
    LUT4 i54005_4_lut (.A(n70763), .B(n23577), .C(n70762), .D(diffExp[0]), 
         .Z(n66912)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i54005_4_lut.init = 16'h5044;
    LUT4 mux_3878_i23_3_lut (.A(\B_int[22] ), .B(\A_int[22] ), .C(diffExpAB[8]), 
         .Z(efectFracB[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3878_i23_3_lut.init = 16'hcaca;
    LUT4 mux_2994_i5_3_lut (.A(diffExpAB[4]), .B(diffExpBA[4]), .C(diffExpAB[8]), 
         .Z(\diffExp[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2994_i5_3_lut.init = 16'hcaca;
    LUT4 mux_2994_i3_3_lut (.A(diffExpAB[2]), .B(diffExpBA[2]), .C(diffExpAB[8]), 
         .Z(\diffExp[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2994_i3_3_lut.init = 16'hcaca;
    LUT4 mux_2994_i2_3_lut (.A(diffExpAB[1]), .B(diffExpBA[1]), .C(diffExpAB[8]), 
         .Z(\diffExp[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2994_i2_3_lut.init = 16'hcaca;
    LUT4 mux_2994_i1_3_lut (.A(diffExpAB[0]), .B(diffExpBA[0]), .C(diffExpAB[8]), 
         .Z(diffExp[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2994_i1_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(n7), .B(n70734), .C(diffExp[0]), .D(\diffExp[1] ), 
         .Z(n66221)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i23877_3_lut (.A(\A_int[18] ), .B(n458), .C(n70727), .Z(n35487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23877_3_lut.init = 16'hcaca;
    LUT4 i23878_3_lut (.A(\B_int[18] ), .B(n35487), .C(n61), .Z(\frac[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23878_3_lut.init = 16'hcaca;
    LUT4 i23872_3_lut (.A(\A_int[13] ), .B(n463), .C(n70727), .Z(n35482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23872_3_lut.init = 16'hcaca;
    LUT4 i23873_3_lut (.A(\B_int[13] ), .B(n35482), .C(n61), .Z(\frac[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23873_3_lut.init = 16'hcaca;
    PFUMX mux_3928_i16 (.BLUT(n37[15]), .ALUT(n37[19]), .C0(\diffExp[2] ), 
          .Z(n69[15]));
    PFUMX mux_3928_i17 (.BLUT(n37[16]), .ALUT(n37[20]), .C0(\diffExp[2] ), 
          .Z(n69[16]));
    PFUMX mux_3928_i18 (.BLUT(n37[17]), .ALUT(n28), .C0(\diffExp[2] ), 
          .Z(n69[17]));
    PFUMX mux_3928_i19 (.BLUT(n37[18]), .ALUT(n37[22]), .C0(\diffExp[2] ), 
          .Z(n69[18]));
    PFUMX mux_3933_i22 (.BLUT(n69[21]), .ALUT(n69[23]), .C0(\diffExp[1] ), 
          .Z(n101[21]));
    PFUMX mux_3933_i23 (.BLUT(n66597), .ALUT(n69[24]), .C0(\diffExp[1] ), 
          .Z(n101[22]));
    PFUMX i56078 (.BLUT(n70872), .ALUT(n70873), .C0(diffExpAB[8]), .Z(n7));
    LUT4 i3_4_lut_else_4_lut (.A(diffExpAB[5]), .B(diffExpAB[7]), .C(diffExpAB[6]), 
         .Z(n70872)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_4_lut_else_4_lut.init = 16'hfefe;
    LUT4 i3_4_lut_then_4_lut (.A(diffExpBA[7]), .B(diffExpBA[8]), .C(diffExpBA[6]), 
         .D(diffExpBA[5]), .Z(n70873)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_then_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module \fp_mul(32,24,8) 
//

module \fp_mul(32,24,8)  (\B_int[12] , \B_int[13] , \B_int[15] , \B_int[8] , 
            \A_int[2] , \A_int[3] , \A_int[6] , \A_int[7] , \A_int[4] , 
            \A_int[5] , \B_int[0] , clock, n73813, alu_b, \A_int[0] , 
            alu_a, \A_int[11] , \A_int[12] , \A_int[13] , \A_int[15] , 
            \A_int[17] , \A_int[16] , \A_int[18] , \A_int[19] , \A_int[14] , 
            n4, n41520, \A_int[1] , \A_int[10] , \A_int[9] , \A_int[22] , 
            \A_int[21] , \A_int[8] , \A_int[20] , n22310, \B_int[11] , 
            \B_int[14] , \B_int[10] , \B_int[9] , \B_int[19] , \B_int[18] , 
            \B_int[20] , \B_int[21] , \B_int[7] , n22437, \prod[47] , 
            n66955, n67025, n67007, n41808, \prod[45] , \prod[46] , 
            \prod[28] , \prod[33] , \prod[40] , \prod[22] , \prod[24] , 
            \prod[25] , \prod[23] , \prod[26] , \prod[41] , \prod[34] , 
            \prod[37] , \prod[27] , \prod[39] , \prod[29] , \prod[35] , 
            \prod[36] , \prod[31] , \prod[32] , \prod[43] , \prod[30] , 
            \prod[38] , \prod[42] , \prod[44] , n42939, n42941, n25571, 
            n73812, n42934, mul_c, GND_net, \frac_norm[20] , \frac_norm[16] , 
            \frac_norm[14] , \frac_norm[15] , \frac_norm[12] , \frac_norm[13] , 
            \frac_norm[10] , \frac_norm[11] , \frac_norm[8] , n15, \B_int[17] , 
            \B_int[16] , \B_int[22] , \frac_norm[7] , n25583, n984, 
            \B_int[3] , \B_int[1] , \B_int[2] , \frac_norm[4] , \frac_norm[5] , 
            \frac_norm[3] , \frac_norm[2] , exp_final, \FP_Z_int[22] , 
            mul_ce, \B_int[6] , \B_int[5] , \B_int[4] , n6, \prod[21] );
    output \B_int[12] ;
    output \B_int[13] ;
    output \B_int[15] ;
    output \B_int[8] ;
    output \A_int[2] ;
    output \A_int[3] ;
    output \A_int[6] ;
    output \A_int[7] ;
    output \A_int[4] ;
    output \A_int[5] ;
    output \B_int[0] ;
    input clock;
    input n73813;
    input [31:0]alu_b;
    output \A_int[0] ;
    input [31:0]alu_a;
    output \A_int[11] ;
    output \A_int[12] ;
    output \A_int[13] ;
    output \A_int[15] ;
    output \A_int[17] ;
    output \A_int[16] ;
    output \A_int[18] ;
    output \A_int[19] ;
    output \A_int[14] ;
    output n4;
    output n41520;
    output \A_int[1] ;
    output \A_int[10] ;
    output \A_int[9] ;
    output \A_int[22] ;
    output \A_int[21] ;
    output \A_int[8] ;
    output \A_int[20] ;
    output n22310;
    output \B_int[11] ;
    output \B_int[14] ;
    output \B_int[10] ;
    output \B_int[9] ;
    output \B_int[19] ;
    output \B_int[18] ;
    output \B_int[20] ;
    output \B_int[21] ;
    output \B_int[7] ;
    output n22437;
    input \prod[47] ;
    input n66955;
    input n67025;
    input n67007;
    output n41808;
    input \prod[45] ;
    input \prod[46] ;
    input \prod[28] ;
    input \prod[33] ;
    input \prod[40] ;
    input \prod[22] ;
    input \prod[24] ;
    input \prod[25] ;
    input \prod[23] ;
    input \prod[26] ;
    input \prod[41] ;
    input \prod[34] ;
    input \prod[37] ;
    input \prod[27] ;
    input \prod[39] ;
    input \prod[29] ;
    input \prod[35] ;
    input \prod[36] ;
    input \prod[31] ;
    input \prod[32] ;
    input \prod[43] ;
    input \prod[30] ;
    input \prod[38] ;
    input \prod[42] ;
    input \prod[44] ;
    output n42939;
    output n42941;
    output n25571;
    input n73812;
    input n42934;
    output [31:0]mul_c;
    input GND_net;
    input \frac_norm[20] ;
    input \frac_norm[16] ;
    input \frac_norm[14] ;
    input \frac_norm[15] ;
    input \frac_norm[12] ;
    input \frac_norm[13] ;
    input \frac_norm[10] ;
    input \frac_norm[11] ;
    input \frac_norm[8] ;
    input n15;
    output \B_int[17] ;
    output \B_int[16] ;
    output \B_int[22] ;
    input \frac_norm[7] ;
    input n25583;
    input [7:0]n984;
    output \B_int[3] ;
    output \B_int[1] ;
    output \B_int[2] ;
    input \frac_norm[4] ;
    input \frac_norm[5] ;
    input \frac_norm[3] ;
    input \frac_norm[2] ;
    output [7:0]exp_final;
    input \FP_Z_int[22] ;
    input mul_ce;
    output \B_int[6] ;
    output \B_int[5] ;
    output \B_int[4] ;
    output n6;
    input \prod[21] ;
    
    wire [31:0]A_int;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(44[11:16])
    wire [31:0]B_int;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(44[18:23])
    wire [7:0]exp_stg2;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(56[11:19])
    wire [7:0]exp_int;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(56[30:37])
    wire [23:0]frac_round;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(64[11:21])
    wire [26:0]frac_norm;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(63[11:20])
    wire [30:0]\sticky_gen.firstOne_B ;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(116[28:38])
    wire [30:0]\sticky_gen.firstOne_A ;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(116[16:26])
    wire sign_stg2;   // c:/users/yisong/documents/new/mlp/fp_mul.vhd(59[11:20])
    
    wire n66190, n14, n70840, n137, n70839, n66601, n6_c, n70838, 
        n4_c, n57, n254, n70825, n70826, n66991, n66969, n70766, 
        n67010, n66763;
    wire [3:0]n261;
    
    wire n70831, n278, n70829, n70830;
    wire [3:0]n279;
    
    wire n66927, n70827, n62771, n70828, n10, n14_adj_469, n66194, 
        n4_adj_470, n41626, n4_adj_471, n15_c, n62828, n10_adj_473, 
        n14_adj_474, n22, n28, n18, n26, n30, n17, n66722, n66179, 
        n12, n66723, n6_adj_475, n70808, n66187, n14_adj_476, n15_adj_477, 
        n10_adj_478, n14_adj_479, n9, n22435, n66755, n36, n30_adj_480, 
        n29, n37, n41, n40, n31, n44, n43, n26242, n9_adj_481, 
        n14_adj_482, n66191, n24070, n70854, n70852, n61588, n61587, 
        n61586, n61585, n61584, n61583, n61582, n6_adj_483, n70608, 
        n61581, n61580, n70780, n61579, n70741, n67053, n70853, 
        n70143, n23, n70141, n70139;
    wire [2:0]n346;
    
    wire n70765, n70140, n70138, n70137, n70136, n67051, n61578, 
        n64329, n63205, n61577, n61576, n61575, n61574, n61572, 
        n61571, n61570, n70742, n73794, n4_adj_485, n70720;
    wire [4:0]n418;
    
    wire n70711;
    wire [31:0]n65;
    wire [31:0]n65_adj_489;
    
    wire n70702, n70696, n8, n66531, n12_adj_487, n6_adj_488, n25, 
        n97, n39740, n39744, n63126, n16;
    
    LUT4 i5_3_lut_4_lut (.A(A_int[30]), .B(B_int[30]), .C(exp_stg2[5]), 
         .D(n66190), .Z(n14)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i5_3_lut_4_lut.init = 16'he000;
    LUT4 i120_2_lut_rep_870 (.A(A_int[30]), .B(B_int[30]), .Z(n70840)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i120_2_lut_rep_870.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(\B_int[12] ), .B(\B_int[13] ), .C(\B_int[15] ), 
         .D(\B_int[8] ), .Z(n137)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_869 (.A(\B_int[12] ), .B(\B_int[13] ), .Z(n70839)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_869.init = 16'heeee;
    LUT4 i2_2_lut_3_lut (.A(\A_int[2] ), .B(\A_int[3] ), .C(n66601), .Z(n6_c)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_868 (.A(\A_int[2] ), .B(\A_int[3] ), .Z(n70838)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_868.init = 16'heeee;
    LUT4 i2_3_lut_4_lut_adj_845 (.A(\A_int[6] ), .B(\A_int[7] ), .C(\A_int[4] ), 
         .D(\A_int[5] ), .Z(n4_c)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_845.init = 16'h000e;
    LUT4 i2_3_lut_4_lut_adj_846 (.A(\A_int[6] ), .B(\A_int[7] ), .C(\A_int[4] ), 
         .D(\A_int[5] ), .Z(n57)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_846.init = 16'hfffe;
    FD1P3AX B_int_i0_i0 (.D(alu_b[0]), .SP(n73813), .CK(clock), .Q(\B_int[0] ));
    defparam B_int_i0_i0.GSR = "DISABLED";
    FD1P3AX A_int_i0_i0 (.D(alu_a[0]), .SP(n73813), .CK(clock), .Q(\A_int[0] ));
    defparam A_int_i0_i0.GSR = "DISABLED";
    LUT4 i54_2_lut_rep_855_3_lut (.A(n254), .B(\A_int[11] ), .C(\A_int[12] ), 
         .Z(n70825)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i54_2_lut_rep_855_3_lut.init = 16'hfefe;
    LUT4 i56_2_lut_3_lut_rep_856_4_lut (.A(n254), .B(\A_int[11] ), .C(\A_int[13] ), 
         .D(\A_int[12] ), .Z(n70826)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i56_2_lut_3_lut_rep_856_4_lut.init = 16'hfffe;
    PFUMX i23 (.BLUT(n66991), .ALUT(n66969), .C0(n70766), .Z(n67010));
    LUT4 i27761_4_lut_4_lut (.A(n254), .B(\A_int[11] ), .C(n66601), .D(n66763), 
         .Z(n261[0])) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam i27761_4_lut_4_lut.init = 16'he444;
    LUT4 i52_2_lut_rep_861 (.A(n254), .B(\A_int[11] ), .Z(n70831)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i52_2_lut_rep_861.init = 16'heeee;
    LUT4 i64_2_lut_3_lut_rep_859_4_lut (.A(n278), .B(\A_int[15] ), .C(\A_int[17] ), 
         .D(\A_int[16] ), .Z(n70829)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i64_2_lut_3_lut_rep_859_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_1_lut_2_lut (.A(n278), .B(\A_int[15] ), .Z(n70830)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_1_lut_2_lut.init = 16'heeee;
    LUT4 i54019_4_lut_4_lut_4_lut (.A(n70830), .B(\A_int[16] ), .C(\A_int[17] ), 
         .D(n279[0]), .Z(n66927)) /* synthesis lut_function=(A (D)+!A !(B+!(C))) */ ;
    defparam i54019_4_lut_4_lut_4_lut.init = 16'hba10;
    LUT4 i66_2_lut_rep_857_4_lut (.A(n70830), .B(\A_int[16] ), .C(\A_int[17] ), 
         .D(\A_int[18] ), .Z(n70827)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i66_2_lut_rep_857_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n70829), .B(\A_int[18] ), .C(\A_int[19] ), 
         .D(n70830), .Z(n62771)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 i68_2_lut_3_lut_rep_858 (.A(n70829), .B(\A_int[18] ), .C(\A_int[19] ), 
         .Z(n70828)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i68_2_lut_3_lut_rep_858.init = 16'hfefe;
    LUT4 i2_2_lut (.A(B_int[25]), .B(B_int[27]), .Z(n10)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(B_int[26]), .B(B_int[24]), .C(B_int[28]), .D(B_int[30]), 
         .Z(n14_adj_469)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i58_2_lut_4_lut (.A(n70831), .B(\A_int[12] ), .C(\A_int[13] ), 
         .D(\A_int[14] ), .Z(n278)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i58_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_847 (.A(n70831), .B(\A_int[12] ), .C(\A_int[13] ), 
         .D(n66194), .Z(n4_adj_470)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_847.init = 16'hfe00;
    LUT4 i7_4_lut (.A(B_int[23]), .B(n14_adj_469), .C(n10), .D(B_int[29]), 
         .Z(n41626)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(B_int[30]), .B(A_int[30]), .Z(n4_adj_471)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i8_4_lut (.A(n15_c), .B(exp_stg2[6]), .C(n14), .D(exp_stg2[1]), 
         .Z(n62828)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(n62828), .B(n41626), .C(exp_int[7]), .D(n4_adj_471), 
         .Z(n4)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfeee;
    LUT4 i2_2_lut_adj_848 (.A(A_int[25]), .B(A_int[29]), .Z(n10_adj_473)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_848.init = 16'h8888;
    LUT4 i6_4_lut_adj_849 (.A(A_int[28]), .B(A_int[30]), .C(A_int[23]), 
         .D(A_int[27]), .Z(n14_adj_474)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_849.init = 16'h8000;
    LUT4 i7_4_lut_adj_850 (.A(A_int[24]), .B(n14_adj_474), .C(n10_adj_473), 
         .D(A_int[26]), .Z(n41520)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_850.init = 16'h8000;
    LUT4 i3_4_lut (.A(n70838), .B(\A_int[0] ), .C(\A_int[1] ), .D(n57), 
         .Z(n66194)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(\A_int[14] ), .B(\A_int[10] ), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(\A_int[16] ), .B(\A_int[11] ), .C(\A_int[13] ), 
         .D(n66194), .Z(n28)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_adj_851 (.A(\A_int[15] ), .B(\A_int[12] ), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_851.init = 16'heeee;
    LUT4 i10_4_lut (.A(\A_int[19] ), .B(\A_int[9] ), .C(\A_int[22] ), 
         .D(\A_int[17] ), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(\A_int[18] ), .B(n28), .C(n22), .D(\A_int[21] ), 
         .Z(n30)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_852 (.A(\A_int[8] ), .B(\A_int[20] ), .Z(n17)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_852.init = 16'heeee;
    LUT4 i15_4_lut (.A(n17), .B(n30), .C(n26), .D(n18), .Z(n22310)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut (.A(\B_int[11] ), .B(\B_int[14] ), .C(\B_int[10] ), 
         .Z(n66722)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i5_4_lut (.A(\B_int[9] ), .B(\B_int[19] ), .C(\B_int[18] ), .D(n66179), 
         .Z(n12)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut_adj_853 (.A(n66722), .B(n12), .C(\B_int[20] ), .D(\B_int[21] ), 
         .Z(n66723)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_853.init = 16'hfffe;
    LUT4 i3_4_lut_adj_854 (.A(n66723), .B(n6_adj_475), .C(\B_int[7] ), 
         .D(n70808), .Z(n66187)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_854.init = 16'hfffe;
    LUT4 i5_3_lut (.A(n66187), .B(B_int[24]), .C(B_int[23]), .Z(n14_adj_476)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut.init = 16'hfefe;
    LUT4 i6_4_lut_adj_855 (.A(B_int[25]), .B(B_int[30]), .C(B_int[26]), 
         .D(B_int[28]), .Z(n15_adj_477)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_855.init = 16'hfffe;
    LUT4 i8_4_lut_adj_856 (.A(n15_adj_477), .B(B_int[27]), .C(n14_adj_476), 
         .D(B_int[29]), .Z(n22437)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut_adj_856.init = 16'hfffe;
    LUT4 i2_2_lut_adj_857 (.A(A_int[27]), .B(A_int[28]), .Z(n10_adj_478)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_857.init = 16'heeee;
    LUT4 i6_4_lut_adj_858 (.A(A_int[25]), .B(A_int[30]), .C(A_int[24]), 
         .D(A_int[26]), .Z(n14_adj_479)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_858.init = 16'hfffe;
    LUT4 i1_2_lut_adj_859 (.A(A_int[23]), .B(A_int[29]), .Z(n9)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_859.init = 16'heeee;
    LUT4 i1_4_lut_adj_860 (.A(n9), .B(n22310), .C(n14_adj_479), .D(n10_adj_478), 
         .Z(n22435)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_860.init = 16'hfffe;
    LUT4 i1_4_lut_adj_861 (.A(\prod[47] ), .B(n66955), .C(n67025), .D(n67007), 
         .Z(n66755)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_861.init = 16'hfffe;
    LUT4 i2_3_lut_adj_862 (.A(n22435), .B(n22437), .C(n66755), .Z(n41808)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_adj_862.init = 16'h8080;
    LUT4 i13_4_lut (.A(\prod[45] ), .B(\prod[46] ), .C(\prod[28] ), .D(\prod[33] ), 
         .Z(n36)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13_4_lut.init = 16'h8000;
    LUT4 i7_2_lut (.A(\prod[40] ), .B(\prod[22] ), .Z(n30_adj_480)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7_2_lut.init = 16'h8888;
    LUT4 i6_2_lut_adj_863 (.A(\prod[24] ), .B(\prod[25] ), .Z(n29)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6_2_lut_adj_863.init = 16'h8888;
    LUT4 i14_4_lut_adj_864 (.A(\prod[23] ), .B(\prod[26] ), .C(\prod[41] ), 
         .D(\prod[34] ), .Z(n37)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i14_4_lut_adj_864.init = 16'h8000;
    LUT4 i18_4_lut (.A(\prod[37] ), .B(n36), .C(\prod[27] ), .D(\prod[39] ), 
         .Z(n41)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(\prod[29] ), .B(\prod[35] ), .C(\prod[36] ), .D(\prod[31] ), 
         .Z(n40)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17_4_lut.init = 16'h8000;
    LUT4 i8_2_lut (.A(\prod[32] ), .B(\prod[43] ), .Z(n31)) /* synthesis lut_function=(A (B)) */ ;
    defparam i8_2_lut.init = 16'h8888;
    LUT4 i21_4_lut (.A(n41), .B(n37), .C(n29), .D(n30_adj_480), .Z(n44)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21_4_lut.init = 16'h8000;
    LUT4 i20_4_lut (.A(n31), .B(n40), .C(\prod[30] ), .D(\prod[38] ), 
         .Z(n43)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20_4_lut.init = 16'h8000;
    LUT4 i2_4_lut (.A(\prod[42] ), .B(n43), .C(\prod[44] ), .D(n44), 
         .Z(n26242)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'h8000;
    LUT4 i2_4_lut_adj_865 (.A(n26242), .B(\prod[47] ), .C(A_int[23]), 
         .D(B_int[23]), .Z(n66190)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;
    defparam i2_4_lut_adj_865.init = 16'hfeef;
    LUT4 i1_2_lut_adj_866 (.A(exp_stg2[2]), .B(exp_stg2[6]), .Z(n9_adj_481)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_866.init = 16'heeee;
    LUT4 i7_4_lut_adj_867 (.A(n9_adj_481), .B(n14_adj_482), .C(exp_stg2[1]), 
         .D(n66190), .Z(n66191)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_867.init = 16'hfffe;
    LUT4 i1_4_lut_adj_868 (.A(n41808), .B(n66191), .C(exp_int[7]), .D(n70840), 
         .Z(n42939)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_868.init = 16'h8880;
    LUT4 i1_3_lut (.A(n41808), .B(n41520), .C(n4), .Z(n42941)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_3_lut.init = 16'ha8a8;
    LUT4 i1_3_lut_adj_869 (.A(n41626), .B(n22435), .C(n66187), .Z(n25571)) /* synthesis lut_function=(A ((C)+!B)) */ ;
    defparam i1_3_lut_adj_869.init = 16'ha2a2;
    LUT4 i12399_4_lut (.A(n73812), .B(n42934), .C(n42941), .D(n42939), 
         .Z(n24070)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;
    defparam i12399_4_lut.init = 16'ha8aa;
    FD1P3IX FP_Z_i0_i1 (.D(frac_round[1]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[1]));
    defparam FP_Z_i0_i1.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i2 (.D(frac_round[2]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[2]));
    defparam FP_Z_i0_i2.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i3 (.D(frac_round[3]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[3]));
    defparam FP_Z_i0_i3.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i4 (.D(frac_round[4]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[4]));
    defparam FP_Z_i0_i4.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i5 (.D(frac_round[5]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[5]));
    defparam FP_Z_i0_i5.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i6 (.D(frac_round[6]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[6]));
    defparam FP_Z_i0_i6.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i7 (.D(frac_round[7]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[7]));
    defparam FP_Z_i0_i7.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_rep_796_4_lut (.A(n70854), .B(n70852), .C(\B_int[7] ), 
         .D(n66179), .Z(n70766)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_rep_796_4_lut.init = 16'hfffe;
    FD1P3IX FP_Z_i0_i8 (.D(frac_round[8]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[8]));
    defparam FP_Z_i0_i8.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i9 (.D(frac_round[9]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[9]));
    defparam FP_Z_i0_i9.GSR = "DISABLED";
    CCU2D add_256_23 (.A0(frac_norm[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(frac_norm[25]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61588), .S0(frac_round[21]), .S1(frac_round[22]));
    defparam add_256_23.INIT0 = 16'h5aaa;
    defparam add_256_23.INIT1 = 16'h5aaa;
    defparam add_256_23.INJECT1_0 = "NO";
    defparam add_256_23.INJECT1_1 = "NO";
    FD1P3IX FP_Z_i0_i10 (.D(frac_round[10]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[10]));
    defparam FP_Z_i0_i10.GSR = "DISABLED";
    CCU2D add_256_21 (.A0(frac_norm[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(frac_norm[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61587), .COUT(n61588), .S0(frac_round[19]), 
          .S1(frac_round[20]));
    defparam add_256_21.INIT0 = 16'h5aaa;
    defparam add_256_21.INIT1 = 16'h5aaa;
    defparam add_256_21.INJECT1_0 = "NO";
    defparam add_256_21.INJECT1_1 = "NO";
    CCU2D add_256_19 (.A0(\frac_norm[20] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(frac_norm[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61586), .COUT(n61587), .S0(frac_round[17]), 
          .S1(frac_round[18]));
    defparam add_256_19.INIT0 = 16'h5aaa;
    defparam add_256_19.INIT1 = 16'h5aaa;
    defparam add_256_19.INJECT1_0 = "NO";
    defparam add_256_19.INJECT1_1 = "NO";
    CCU2D add_256_17 (.A0(frac_norm[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(frac_norm[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61585), .COUT(n61586), .S0(frac_round[15]), 
          .S1(frac_round[16]));
    defparam add_256_17.INIT0 = 16'h5aaa;
    defparam add_256_17.INIT1 = 16'h5aaa;
    defparam add_256_17.INJECT1_0 = "NO";
    defparam add_256_17.INJECT1_1 = "NO";
    CCU2D add_256_15 (.A0(\frac_norm[16] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(frac_norm[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61584), .COUT(n61585), .S0(frac_round[13]), 
          .S1(frac_round[14]));
    defparam add_256_15.INIT0 = 16'h5aaa;
    defparam add_256_15.INIT1 = 16'h5aaa;
    defparam add_256_15.INJECT1_0 = "NO";
    defparam add_256_15.INJECT1_1 = "NO";
    CCU2D add_256_13 (.A0(\frac_norm[14] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\frac_norm[15] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61583), .COUT(n61584), .S0(frac_round[11]), 
          .S1(frac_round[12]));
    defparam add_256_13.INIT0 = 16'h5aaa;
    defparam add_256_13.INIT1 = 16'h5aaa;
    defparam add_256_13.INJECT1_0 = "NO";
    defparam add_256_13.INJECT1_1 = "NO";
    FD1P3IX FP_Z_i0_i11 (.D(frac_round[11]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[11]));
    defparam FP_Z_i0_i11.GSR = "DISABLED";
    CCU2D add_256_11 (.A0(\frac_norm[12] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\frac_norm[13] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61582), .COUT(n61583), .S0(frac_round[9]), 
          .S1(frac_round[10]));
    defparam add_256_11.INIT0 = 16'h5aaa;
    defparam add_256_11.INIT1 = 16'h5aaa;
    defparam add_256_11.INJECT1_0 = "NO";
    defparam add_256_11.INJECT1_1 = "NO";
    LUT4 \sticky_gen.firstOne_B_0__bdd_4_lut  (.A(\sticky_gen.firstOne_B [0]), 
         .B(\sticky_gen.firstOne_B [1]), .C(\sticky_gen.firstOne_A [1]), 
         .D(n6_adj_483), .Z(n70608)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C (D))+!B !(C+!(D)))) */ ;
    defparam \sticky_gen.firstOne_B_0__bdd_4_lut .init = 16'hbed7;
    CCU2D add_256_9 (.A0(\frac_norm[10] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\frac_norm[11] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61581), .COUT(n61582), .S0(frac_round[7]), 
          .S1(frac_round[8]));
    defparam add_256_9.INIT0 = 16'h5aaa;
    defparam add_256_9.INIT1 = 16'h5aaa;
    defparam add_256_9.INJECT1_0 = "NO";
    defparam add_256_9.INJECT1_1 = "NO";
    FD1P3IX FP_Z_i0_i12 (.D(frac_round[12]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[12]));
    defparam FP_Z_i0_i12.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i13 (.D(frac_round[13]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[13]));
    defparam FP_Z_i0_i13.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i14 (.D(frac_round[14]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[14]));
    defparam FP_Z_i0_i14.GSR = "DISABLED";
    CCU2D add_256_7 (.A0(\frac_norm[8] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\prod[30] ), .B1(\prod[47] ), .C1(\prod[29] ), 
          .D1(n15), .CIN(n61580), .COUT(n61581), .S0(frac_round[5]), 
          .S1(frac_round[6]));
    defparam add_256_7.INIT0 = 16'h5aaa;
    defparam add_256_7.INIT1 = 16'hf888;
    defparam add_256_7.INJECT1_0 = "NO";
    defparam add_256_7.INJECT1_1 = "NO";
    LUT4 i6_4_lut_4_lut (.A(exp_int[7]), .B(exp_stg2[3]), .C(exp_stg2[5]), 
         .D(exp_stg2[4]), .Z(n14_adj_482)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i6_4_lut_4_lut.init = 16'hfffd;
    LUT4 i2_2_lut_4_lut (.A(\B_int[17] ), .B(\B_int[16] ), .C(n137), .D(\B_int[22] ), 
         .Z(n6_adj_475)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_rep_810 (.A(\B_int[17] ), .B(\B_int[16] ), .C(n137), 
         .Z(n70780)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_810.init = 16'hfefe;
    FD1P3IX FP_Z_i0_i15 (.D(frac_round[15]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[15]));
    defparam FP_Z_i0_i15.GSR = "DISABLED";
    LUT4 i6_4_lut_4_lut_adj_870 (.A(exp_int[7]), .B(exp_stg2[3]), .C(exp_stg2[4]), 
         .D(exp_stg2[2]), .Z(n15_c)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i6_4_lut_4_lut_adj_870.init = 16'h4000;
    CCU2D add_256_5 (.A0(\prod[27] ), .B0(\prod[47] ), .C0(\prod[26] ), 
          .D0(n15), .A1(\frac_norm[7] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61579), .COUT(n61580), .S0(frac_round[3]), 
          .S1(frac_round[4]));
    defparam add_256_5.INIT0 = 16'hf888;
    defparam add_256_5.INIT1 = 16'h5aaa;
    defparam add_256_5.INJECT1_0 = "NO";
    defparam add_256_5.INJECT1_1 = "NO";
    FD1P3IX FP_Z_i0_i16 (.D(frac_round[16]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[16]));
    defparam FP_Z_i0_i16.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i17 (.D(frac_round[17]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[17]));
    defparam FP_Z_i0_i17.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i18 (.D(frac_round[18]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[18]));
    defparam FP_Z_i0_i18.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i19 (.D(frac_round[19]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[19]));
    defparam FP_Z_i0_i19.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i20 (.D(frac_round[20]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[20]));
    defparam FP_Z_i0_i20.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i21 (.D(frac_round[21]), .SP(n73813), .CD(n24070), 
            .CK(clock), .Q(mul_c[21]));
    defparam FP_Z_i0_i21.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_771_4_lut (.A(n66179), .B(n70808), .C(\B_int[7] ), 
         .D(\B_int[9] ), .Z(n70741)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_771_4_lut.init = 16'hfffe;
    FD1P3JX FP_Z_i0_i23 (.D(n984[0]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[23]));
    defparam FP_Z_i0_i23.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i24 (.D(n984[1]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[24]));
    defparam FP_Z_i0_i24.GSR = "DISABLED";
    LUT4 n67053_bdd_4_lut_56996 (.A(n67053), .B(n70853), .C(\B_int[9] ), 
         .D(\B_int[8] ), .Z(n70143)) /* synthesis lut_function=(!(A (C+(D))+!A ((C)+!B))) */ ;
    defparam n67053_bdd_4_lut_56996.init = 16'h040e;
    LUT4 n23_bdd_4_lut_56073 (.A(n23), .B(\B_int[3] ), .C(\B_int[1] ), 
         .D(\B_int[2] ), .Z(n70141)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam n23_bdd_4_lut_56073.init = 16'h0f0d;
    PFUMX i55881 (.BLUT(n70139), .ALUT(n346[0]), .C0(n70765), .Z(n70140));
    LUT4 n70138_bdd_2_lut_57055 (.A(n70138), .B(\B_int[7] ), .Z(n70139)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n70138_bdd_2_lut_57055.init = 16'heeee;
    PFUMX i55879 (.BLUT(n70137), .ALUT(n70136), .C0(n67051), .Z(n70138));
    LUT4 n67051_bdd_3_lut_56061 (.A(\B_int[10] ), .B(\B_int[11] ), .C(\B_int[9] ), 
         .Z(n70137)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;
    defparam n67051_bdd_3_lut_56061.init = 16'hf4f4;
    LUT4 n67051_bdd_3_lut_55878 (.A(\B_int[10] ), .B(\B_int[9] ), .C(\B_int[8] ), 
         .Z(n70136)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;
    defparam n67051_bdd_3_lut_55878.init = 16'h0d0d;
    FD1P3JX FP_Z_i0_i25 (.D(n984[2]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[25]));
    defparam FP_Z_i0_i25.GSR = "DISABLED";
    CCU2D add_256_3 (.A0(\frac_norm[4] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\frac_norm[5] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61578), .COUT(n61579), .S0(frac_round[1]), 
          .S1(frac_round[2]));
    defparam add_256_3.INIT0 = 16'h5aaa;
    defparam add_256_3.INIT1 = 16'h5aaa;
    defparam add_256_3.INJECT1_0 = "NO";
    defparam add_256_3.INJECT1_1 = "NO";
    CCU2D add_256_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\frac_norm[3] ), .B1(n64329), .C1(n63205), .D1(\frac_norm[2] ), 
          .COUT(n61578), .S1(frac_round[0]));
    defparam add_256_1.INIT0 = 16'hF000;
    defparam add_256_1.INIT1 = 16'h56a6;
    defparam add_256_1.INJECT1_0 = "NO";
    defparam add_256_1.INJECT1_1 = "NO";
    FD1P3JX FP_Z_i0_i26 (.D(n984[3]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[26]));
    defparam FP_Z_i0_i26.GSR = "DISABLED";
    CCU2D add_130_9 (.A0(exp_int[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61577), 
          .S0(exp_final[7]));
    defparam add_130_9.INIT0 = 16'ha555;
    defparam add_130_9.INIT1 = 16'h0000;
    defparam add_130_9.INJECT1_0 = "NO";
    defparam add_130_9.INJECT1_1 = "NO";
    CCU2D add_130_7 (.A0(exp_stg2[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_stg2[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61576), .COUT(n61577), .S0(exp_final[5]), .S1(exp_final[6]));
    defparam add_130_7.INIT0 = 16'h5aaa;
    defparam add_130_7.INIT1 = 16'h5aaa;
    defparam add_130_7.INJECT1_0 = "NO";
    defparam add_130_7.INJECT1_1 = "NO";
    FD1P3JX FP_Z_i0_i27 (.D(n984[4]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[27]));
    defparam FP_Z_i0_i27.GSR = "DISABLED";
    CCU2D add_130_5 (.A0(exp_stg2[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_stg2[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61575), .COUT(n61576), .S0(exp_final[3]), .S1(exp_final[4]));
    defparam add_130_5.INIT0 = 16'h5aaa;
    defparam add_130_5.INIT1 = 16'h5aaa;
    defparam add_130_5.INJECT1_0 = "NO";
    defparam add_130_5.INJECT1_1 = "NO";
    FD1P3JX FP_Z_i0_i28 (.D(n984[5]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[28]));
    defparam FP_Z_i0_i28.GSR = "DISABLED";
    CCU2D add_130_3 (.A0(exp_stg2[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_stg2[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61574), .COUT(n61575), .S0(exp_final[1]), .S1(exp_final[2]));
    defparam add_130_3.INIT0 = 16'h5aaa;
    defparam add_130_3.INIT1 = 16'h5aaa;
    defparam add_130_3.INJECT1_0 = "NO";
    defparam add_130_3.INJECT1_1 = "NO";
    CCU2D add_130_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[23]), .B1(B_int[23]), .C1(n26242), .D1(\prod[47] ), 
          .COUT(n61574), .S1(exp_final[0]));
    defparam add_130_1.INIT0 = 16'hF000;
    defparam add_130_1.INIT1 = 16'h6669;
    defparam add_130_1.INJECT1_0 = "NO";
    defparam add_130_1.INJECT1_1 = "NO";
    FD1P3JX FP_Z_i0_i29 (.D(n984[6]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[29]));
    defparam FP_Z_i0_i29.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i30 (.D(n984[7]), .SP(n73813), .PD(n25583), .CK(clock), 
            .Q(mul_c[30]));
    defparam FP_Z_i0_i30.GSR = "DISABLED";
    CCU2D add_114_8 (.A0(A_int[29]), .B0(B_int[29]), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[30]), .B1(B_int[30]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61572), .S0(exp_stg2[6]), .S1(exp_int[7]));
    defparam add_114_8.INIT0 = 16'h5666;
    defparam add_114_8.INIT1 = 16'h5666;
    defparam add_114_8.INJECT1_0 = "NO";
    defparam add_114_8.INJECT1_1 = "NO";
    CCU2D add_114_6 (.A0(A_int[27]), .B0(B_int[27]), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[28]), .B1(B_int[28]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61571), .COUT(n61572), .S0(exp_stg2[4]), .S1(exp_stg2[5]));
    defparam add_114_6.INIT0 = 16'h5666;
    defparam add_114_6.INIT1 = 16'h5666;
    defparam add_114_6.INJECT1_0 = "NO";
    defparam add_114_6.INJECT1_1 = "NO";
    CCU2D add_114_4 (.A0(A_int[25]), .B0(B_int[25]), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[26]), .B1(B_int[26]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61570), .COUT(n61571), .S0(exp_stg2[2]), .S1(exp_stg2[3]));
    defparam add_114_4.INIT0 = 16'h5666;
    defparam add_114_4.INIT1 = 16'h5666;
    defparam add_114_4.INJECT1_0 = "NO";
    defparam add_114_4.INJECT1_1 = "NO";
    CCU2D add_114_2 (.A0(A_int[23]), .B0(B_int[23]), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[24]), .B1(B_int[24]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61570), .S1(exp_stg2[1]));
    defparam add_114_2.INIT0 = 16'h1000;
    defparam add_114_2.INIT1 = 16'h5666;
    defparam add_114_2.INJECT1_0 = "NO";
    defparam add_114_2.INJECT1_1 = "NO";
    LUT4 i50_2_lut_4_lut (.A(\A_int[8] ), .B(\A_int[9] ), .C(n66194), 
         .D(\A_int[10] ), .Z(n254)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i50_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_871 (.A(\A_int[8] ), .B(\A_int[9] ), .C(n66194), 
         .D(\A_int[0] ), .Z(n66601)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i1_2_lut_4_lut_adj_871.init = 16'h00fe;
    LUT4 i48_3_lut_rep_772 (.A(\A_int[8] ), .B(\A_int[9] ), .C(n66194), 
         .Z(n70742)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i48_3_lut_rep_772.init = 16'hfefe;
    LUT4 n70141_bdd_4_lut (.A(n70141), .B(\B_int[0] ), .C(n70143), .D(n70766), 
         .Z(n73794)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n70141_bdd_4_lut.init = 16'h22f0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\B_int[9] ), .B(n70766), .C(n137), .D(n66722), 
         .Z(n4_adj_485)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_750_3_lut_4_lut (.A(\B_int[9] ), .B(n70766), .C(n70780), 
         .D(n66722), .Z(n70720)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_750_3_lut_4_lut.init = 16'hfffe;
    FD1P3AX FP_Z_i0_i31 (.D(sign_stg2), .SP(n73813), .CK(clock), .Q(mul_c[31]));
    defparam FP_Z_i0_i31.GSR = "DISABLED";
    FD1P3AX FP_Z_i0_i22 (.D(\FP_Z_int[22] ), .SP(n73813), .CK(clock), 
            .Q(mul_c[22]));
    defparam FP_Z_i0_i22.GSR = "DISABLED";
    FD1P3AX A_int_i0_i30 (.D(alu_a[30]), .SP(n73813), .CK(clock), .Q(A_int[30]));
    defparam A_int_i0_i30.GSR = "DISABLED";
    FD1P3AX A_int_i0_i29 (.D(alu_a[29]), .SP(n73813), .CK(clock), .Q(A_int[29]));
    defparam A_int_i0_i29.GSR = "DISABLED";
    FD1P3AX A_int_i0_i28 (.D(alu_a[28]), .SP(n73813), .CK(clock), .Q(A_int[28]));
    defparam A_int_i0_i28.GSR = "DISABLED";
    FD1P3AX A_int_i0_i27 (.D(alu_a[27]), .SP(n73813), .CK(clock), .Q(A_int[27]));
    defparam A_int_i0_i27.GSR = "DISABLED";
    FD1P3AX A_int_i0_i26 (.D(alu_a[26]), .SP(n73813), .CK(clock), .Q(A_int[26]));
    defparam A_int_i0_i26.GSR = "DISABLED";
    FD1P3AX A_int_i0_i25 (.D(alu_a[25]), .SP(n73813), .CK(clock), .Q(A_int[25]));
    defparam A_int_i0_i25.GSR = "DISABLED";
    FD1P3AX A_int_i0_i24 (.D(alu_a[24]), .SP(n73813), .CK(clock), .Q(A_int[24]));
    defparam A_int_i0_i24.GSR = "DISABLED";
    FD1P3AX A_int_i0_i23 (.D(alu_a[23]), .SP(n73813), .CK(clock), .Q(A_int[23]));
    defparam A_int_i0_i23.GSR = "DISABLED";
    FD1P3AX A_int_i0_i22 (.D(alu_a[22]), .SP(n73813), .CK(clock), .Q(\A_int[22] ));
    defparam A_int_i0_i22.GSR = "DISABLED";
    FD1P3AX A_int_i0_i21 (.D(alu_a[21]), .SP(n73813), .CK(clock), .Q(\A_int[21] ));
    defparam A_int_i0_i21.GSR = "DISABLED";
    FD1P3AX A_int_i0_i20 (.D(alu_a[20]), .SP(n73813), .CK(clock), .Q(\A_int[20] ));
    defparam A_int_i0_i20.GSR = "DISABLED";
    FD1P3AX A_int_i0_i19 (.D(alu_a[19]), .SP(n73813), .CK(clock), .Q(\A_int[19] ));
    defparam A_int_i0_i19.GSR = "DISABLED";
    FD1P3AX A_int_i0_i18 (.D(alu_a[18]), .SP(n73813), .CK(clock), .Q(\A_int[18] ));
    defparam A_int_i0_i18.GSR = "DISABLED";
    FD1P3AX A_int_i0_i17 (.D(alu_a[17]), .SP(n73813), .CK(clock), .Q(\A_int[17] ));
    defparam A_int_i0_i17.GSR = "DISABLED";
    FD1P3AX A_int_i0_i16 (.D(alu_a[16]), .SP(n73813), .CK(clock), .Q(\A_int[16] ));
    defparam A_int_i0_i16.GSR = "DISABLED";
    FD1P3AX A_int_i0_i15 (.D(alu_a[15]), .SP(n73813), .CK(clock), .Q(\A_int[15] ));
    defparam A_int_i0_i15.GSR = "DISABLED";
    FD1P3AX A_int_i0_i14 (.D(alu_a[14]), .SP(mul_ce), .CK(clock), .Q(\A_int[14] ));
    defparam A_int_i0_i14.GSR = "DISABLED";
    FD1P3AX A_int_i0_i13 (.D(alu_a[13]), .SP(mul_ce), .CK(clock), .Q(\A_int[13] ));
    defparam A_int_i0_i13.GSR = "DISABLED";
    FD1P3AX A_int_i0_i12 (.D(alu_a[12]), .SP(mul_ce), .CK(clock), .Q(\A_int[12] ));
    defparam A_int_i0_i12.GSR = "DISABLED";
    FD1P3AX A_int_i0_i11 (.D(alu_a[11]), .SP(mul_ce), .CK(clock), .Q(\A_int[11] ));
    defparam A_int_i0_i11.GSR = "DISABLED";
    FD1P3AX A_int_i0_i10 (.D(alu_a[10]), .SP(mul_ce), .CK(clock), .Q(\A_int[10] ));
    defparam A_int_i0_i10.GSR = "DISABLED";
    FD1P3AX A_int_i0_i9 (.D(alu_a[9]), .SP(mul_ce), .CK(clock), .Q(\A_int[9] ));
    defparam A_int_i0_i9.GSR = "DISABLED";
    FD1P3AX A_int_i0_i8 (.D(alu_a[8]), .SP(mul_ce), .CK(clock), .Q(\A_int[8] ));
    defparam A_int_i0_i8.GSR = "DISABLED";
    FD1P3AX A_int_i0_i7 (.D(alu_a[7]), .SP(mul_ce), .CK(clock), .Q(\A_int[7] ));
    defparam A_int_i0_i7.GSR = "DISABLED";
    FD1P3AX A_int_i0_i6 (.D(alu_a[6]), .SP(mul_ce), .CK(clock), .Q(\A_int[6] ));
    defparam A_int_i0_i6.GSR = "DISABLED";
    FD1P3AX A_int_i0_i5 (.D(alu_a[5]), .SP(mul_ce), .CK(clock), .Q(\A_int[5] ));
    defparam A_int_i0_i5.GSR = "DISABLED";
    FD1P3AX A_int_i0_i4 (.D(alu_a[4]), .SP(mul_ce), .CK(clock), .Q(\A_int[4] ));
    defparam A_int_i0_i4.GSR = "DISABLED";
    FD1P3AX A_int_i0_i3 (.D(alu_a[3]), .SP(mul_ce), .CK(clock), .Q(\A_int[3] ));
    defparam A_int_i0_i3.GSR = "DISABLED";
    FD1P3AX A_int_i0_i2 (.D(alu_a[2]), .SP(mul_ce), .CK(clock), .Q(\A_int[2] ));
    defparam A_int_i0_i2.GSR = "DISABLED";
    FD1P3AX A_int_i0_i1 (.D(alu_a[1]), .SP(mul_ce), .CK(clock), .Q(\A_int[1] ));
    defparam A_int_i0_i1.GSR = "DISABLED";
    FD1P3AX B_int_i0_i30 (.D(alu_b[30]), .SP(mul_ce), .CK(clock), .Q(B_int[30]));
    defparam B_int_i0_i30.GSR = "DISABLED";
    FD1P3AX B_int_i0_i29 (.D(alu_b[29]), .SP(mul_ce), .CK(clock), .Q(B_int[29]));
    defparam B_int_i0_i29.GSR = "DISABLED";
    FD1P3AX B_int_i0_i28 (.D(alu_b[28]), .SP(mul_ce), .CK(clock), .Q(B_int[28]));
    defparam B_int_i0_i28.GSR = "DISABLED";
    FD1P3AX B_int_i0_i27 (.D(alu_b[27]), .SP(mul_ce), .CK(clock), .Q(B_int[27]));
    defparam B_int_i0_i27.GSR = "DISABLED";
    FD1P3AX B_int_i0_i26 (.D(alu_b[26]), .SP(mul_ce), .CK(clock), .Q(B_int[26]));
    defparam B_int_i0_i26.GSR = "DISABLED";
    FD1P3AX B_int_i0_i25 (.D(alu_b[25]), .SP(mul_ce), .CK(clock), .Q(B_int[25]));
    defparam B_int_i0_i25.GSR = "DISABLED";
    FD1P3AX B_int_i0_i24 (.D(alu_b[24]), .SP(mul_ce), .CK(clock), .Q(B_int[24]));
    defparam B_int_i0_i24.GSR = "DISABLED";
    FD1P3AX B_int_i0_i23 (.D(alu_b[23]), .SP(mul_ce), .CK(clock), .Q(B_int[23]));
    defparam B_int_i0_i23.GSR = "DISABLED";
    FD1P3AX B_int_i0_i22 (.D(alu_b[22]), .SP(mul_ce), .CK(clock), .Q(\B_int[22] ));
    defparam B_int_i0_i22.GSR = "DISABLED";
    FD1P3AX B_int_i0_i21 (.D(alu_b[21]), .SP(mul_ce), .CK(clock), .Q(\B_int[21] ));
    defparam B_int_i0_i21.GSR = "DISABLED";
    FD1P3AX B_int_i0_i20 (.D(alu_b[20]), .SP(mul_ce), .CK(clock), .Q(\B_int[20] ));
    defparam B_int_i0_i20.GSR = "DISABLED";
    FD1P3AX B_int_i0_i19 (.D(alu_b[19]), .SP(mul_ce), .CK(clock), .Q(\B_int[19] ));
    defparam B_int_i0_i19.GSR = "DISABLED";
    FD1P3AX B_int_i0_i18 (.D(alu_b[18]), .SP(mul_ce), .CK(clock), .Q(\B_int[18] ));
    defparam B_int_i0_i18.GSR = "DISABLED";
    FD1P3AX B_int_i0_i17 (.D(alu_b[17]), .SP(mul_ce), .CK(clock), .Q(\B_int[17] ));
    defparam B_int_i0_i17.GSR = "DISABLED";
    FD1P3AX B_int_i0_i16 (.D(alu_b[16]), .SP(mul_ce), .CK(clock), .Q(\B_int[16] ));
    defparam B_int_i0_i16.GSR = "DISABLED";
    FD1P3AX B_int_i0_i15 (.D(alu_b[15]), .SP(mul_ce), .CK(clock), .Q(\B_int[15] ));
    defparam B_int_i0_i15.GSR = "DISABLED";
    FD1P3AX B_int_i0_i14 (.D(alu_b[14]), .SP(mul_ce), .CK(clock), .Q(\B_int[14] ));
    defparam B_int_i0_i14.GSR = "DISABLED";
    FD1P3AX B_int_i0_i13 (.D(alu_b[13]), .SP(mul_ce), .CK(clock), .Q(\B_int[13] ));
    defparam B_int_i0_i13.GSR = "DISABLED";
    FD1P3AX B_int_i0_i12 (.D(alu_b[12]), .SP(mul_ce), .CK(clock), .Q(\B_int[12] ));
    defparam B_int_i0_i12.GSR = "DISABLED";
    FD1P3AX B_int_i0_i11 (.D(alu_b[11]), .SP(mul_ce), .CK(clock), .Q(\B_int[11] ));
    defparam B_int_i0_i11.GSR = "DISABLED";
    FD1P3AX B_int_i0_i10 (.D(alu_b[10]), .SP(mul_ce), .CK(clock), .Q(\B_int[10] ));
    defparam B_int_i0_i10.GSR = "DISABLED";
    FD1P3AX B_int_i0_i9 (.D(alu_b[9]), .SP(mul_ce), .CK(clock), .Q(\B_int[9] ));
    defparam B_int_i0_i9.GSR = "DISABLED";
    FD1P3AX B_int_i0_i8 (.D(alu_b[8]), .SP(mul_ce), .CK(clock), .Q(\B_int[8] ));
    defparam B_int_i0_i8.GSR = "DISABLED";
    FD1P3AX B_int_i0_i7 (.D(alu_b[7]), .SP(mul_ce), .CK(clock), .Q(\B_int[7] ));
    defparam B_int_i0_i7.GSR = "DISABLED";
    FD1P3AX B_int_i0_i6 (.D(alu_b[6]), .SP(mul_ce), .CK(clock), .Q(\B_int[6] ));
    defparam B_int_i0_i6.GSR = "DISABLED";
    FD1P3AX B_int_i0_i5 (.D(alu_b[5]), .SP(mul_ce), .CK(clock), .Q(\B_int[5] ));
    defparam B_int_i0_i5.GSR = "DISABLED";
    FD1P3AX B_int_i0_i4 (.D(alu_b[4]), .SP(mul_ce), .CK(clock), .Q(\B_int[4] ));
    defparam B_int_i0_i4.GSR = "DISABLED";
    FD1P3AX B_int_i0_i3 (.D(alu_b[3]), .SP(mul_ce), .CK(clock), .Q(\B_int[3] ));
    defparam B_int_i0_i3.GSR = "DISABLED";
    FD1P3AX B_int_i0_i2 (.D(alu_b[2]), .SP(mul_ce), .CK(clock), .Q(\B_int[2] ));
    defparam B_int_i0_i2.GSR = "DISABLED";
    FD1P3AX B_int_i0_i1 (.D(alu_b[1]), .SP(mul_ce), .CK(clock), .Q(\B_int[1] ));
    defparam B_int_i0_i1.GSR = "DISABLED";
    LUT4 i27776_2_lut_3_lut_4_lut (.A(n70741), .B(n66722), .C(n70140), 
         .D(n70780), .Z(n418[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i27776_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_741_3_lut_4_lut (.A(n70741), .B(n66722), .C(\B_int[18] ), 
         .D(n70780), .Z(n70711)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_741_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_adj_872 (.A(\B_int[6] ), .B(\B_int[0] ), .C(\B_int[5] ), 
         .Z(n66179)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_adj_872.init = 16'hfefe;
    LUT4 i29430_3_lut_4_lut_4_lut (.A(n70720), .B(n73794), .C(n70711), 
         .D(\B_int[19] ), .Z(\sticky_gen.firstOne_B [1])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;
    defparam i29430_3_lut_4_lut_4_lut.init = 16'hddd0;
    LUT4 i2_3_lut_4_lut_adj_873 (.A(\B_int[19] ), .B(n70711), .C(n70766), 
         .D(n4_adj_485), .Z(\sticky_gen.firstOne_B [3])) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut_adj_873.init = 16'h0e00;
    LUT4 i18081_4_lut_4_lut (.A(\B_int[19] ), .B(n70711), .C(n418[0]), 
         .D(\B_int[20] ), .Z(\sticky_gen.firstOne_B [0])) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(D))) */ ;
    defparam i18081_4_lut_4_lut.init = 16'he2f3;
    FD1P3AX B_int_rep_2__i31 (.D(alu_b[31]), .SP(mul_ce), .CK(clock), 
            .Q(n65[31]));
    defparam B_int_rep_2__i31.GSR = "DISABLED";
    LUT4 i29429_3_lut_4_lut (.A(\B_int[19] ), .B(n70711), .C(n67010), 
         .D(n4_adj_485), .Z(\sticky_gen.firstOne_B [2])) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;
    defparam i29429_3_lut_4_lut.init = 16'hf111;
    FD1P3AX A_int_rep_1__i31 (.D(alu_a[31]), .SP(mul_ce), .CK(clock), 
            .Q(n65_adj_489[31]));
    defparam A_int_rep_1__i31.GSR = "DISABLED";
    LUT4 i4925_4_lut_3_lut_rep_732_4_lut (.A(n6_adj_483), .B(\sticky_gen.firstOne_B [0]), 
         .C(\sticky_gen.firstOne_A [1]), .D(\sticky_gen.firstOne_B [1]), 
         .Z(n70702)) /* synthesis lut_function=(A (C (D))+!A (B (C+(D))+!B (C (D)))) */ ;
    defparam i4925_4_lut_3_lut_rep_732_4_lut.init = 16'hf440;
    FD1P3IX FP_Z_i0_i0 (.D(frac_round[0]), .SP(n73813), .CD(n24070), .CK(clock), 
            .Q(mul_c[0]));
    defparam FP_Z_i0_i0.GSR = "DISABLED";
    LUT4 i4932_4_lut_3_lut_rep_726 (.A(\sticky_gen.firstOne_B [2]), .B(n70702), 
         .C(\sticky_gen.firstOne_A [2]), .Z(n70696)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;
    defparam i4932_4_lut_3_lut_rep_726.init = 16'he8e8;
    LUT4 i4939_4_lut_3_lut (.A(\sticky_gen.firstOne_B [3]), .B(n70696), 
         .C(\sticky_gen.firstOne_A [3]), .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;
    defparam i4939_4_lut_3_lut.init = 16'he8e8;
    LUT4 i2_2_lut_adj_874 (.A(frac_round[22]), .B(n41520), .Z(n6)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i2_2_lut_adj_874.init = 16'h2222;
    LUT4 i118_2_lut (.A(n65_adj_489[31]), .B(n65[31]), .Z(sign_stg2)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i118_2_lut.init = 16'h6666;
    LUT4 i2_4_lut_adj_875 (.A(n70830), .B(n70831), .C(n70828), .D(n4_adj_470), 
         .Z(\sticky_gen.firstOne_A [3])) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i2_4_lut_adj_875.init = 16'h20a0;
    LUT4 i55065_3_lut_4_lut (.A(\B_int[1] ), .B(\B_int[3] ), .C(\B_int[2] ), 
         .D(\B_int[0] ), .Z(n66969)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i55065_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_876 (.A(\A_int[1] ), .B(n70831), .C(n6_c), .D(n57), 
         .Z(n66531)) /* synthesis lut_function=(!(A (B)+!A !((C (D))+!B))) */ ;
    defparam i1_4_lut_adj_876.init = 16'h7333;
    LUT4 i29438_4_lut (.A(n70826), .B(n70828), .C(n70830), .D(n66531), 
         .Z(\sticky_gen.firstOne_A [2])) /* synthesis lut_function=(A ((C (D))+!B)+!A ((C)+!B)) */ ;
    defparam i29438_4_lut.init = 16'hf373;
    LUT4 i1_2_lut_rep_838_3_lut_4_lut (.A(\B_int[1] ), .B(\B_int[3] ), .C(\B_int[4] ), 
         .D(\B_int[2] ), .Z(n70808)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_838_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_884 (.A(\B_int[1] ), .B(\B_int[3] ), .Z(n70854)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_884.init = 16'heeee;
    LUT4 i55068_3_lut_4_lut (.A(\B_int[10] ), .B(\B_int[11] ), .C(\B_int[8] ), 
         .D(\B_int[9] ), .Z(n66991)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i55068_3_lut_4_lut.init = 16'h0001;
    LUT4 i53972_2_lut_rep_883 (.A(\B_int[10] ), .B(\B_int[11] ), .Z(n70853)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53972_2_lut_rep_883.init = 16'heeee;
    LUT4 i18075_4_lut_4_lut (.A(\B_int[2] ), .B(\B_int[4] ), .C(\B_int[3] ), 
         .D(\B_int[5] ), .Z(n12_adj_487)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;
    defparam i18075_4_lut_4_lut.init = 16'h5150;
    LUT4 i1_2_lut_adj_877 (.A(\A_int[8] ), .B(\A_int[7] ), .Z(n6_adj_488)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_877.init = 16'h2222;
    LUT4 i1_4_lut_adj_878 (.A(\A_int[4] ), .B(\A_int[5] ), .C(n6_adj_488), 
         .D(\A_int[6] ), .Z(n25)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_878.init = 16'hbbba;
    LUT4 i1_2_lut_rep_795_3_lut_4_lut (.A(\B_int[2] ), .B(\B_int[4] ), .C(n66179), 
         .D(n70854), .Z(n70765)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_795_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_879 (.A(\A_int[1] ), .B(\A_int[2] ), .C(\A_int[3] ), 
         .D(n25), .Z(n66763)) /* synthesis lut_function=(A+!(B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_879.init = 16'hbabb;
    LUT4 i27766_4_lut (.A(n261[0]), .B(n278), .C(n70826), .D(n70825), 
         .Z(n279[0])) /* synthesis lut_function=(A ((C)+!B)+!A !(B ((D)+!C))) */ ;
    defparam i27766_4_lut.init = 16'hb3f3;
    LUT4 i1_2_lut_rep_882 (.A(\B_int[2] ), .B(\B_int[4] ), .Z(n70852)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_882.init = 16'heeee;
    LUT4 i14_4_lut_adj_880 (.A(\A_int[20] ), .B(n66927), .C(n70828), .D(n70827), 
         .Z(n6_adj_483)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i14_4_lut_adj_880.init = 16'h3a0a;
    LUT4 i1_4_lut_adj_881 (.A(\A_int[0] ), .B(\A_int[1] ), .C(n4_c), .D(n70838), 
         .Z(n97)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_881.init = 16'heeef;
    LUT4 i29448_4_lut (.A(n70742), .B(n70826), .C(n70831), .D(n97), 
         .Z(n279[1])) /* synthesis lut_function=(!(A (B ((D)+!C))+!A !((C)+!B))) */ ;
    defparam i29448_4_lut.init = 16'h73f3;
    LUT4 i29439_4_lut (.A(n279[1]), .B(n70828), .C(n70829), .D(n70830), 
         .Z(\sticky_gen.firstOne_A [1])) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;
    defparam i29439_4_lut.init = 16'h8c0c;
    LUT4 i28147_4_lut (.A(n70608), .B(n70702), .C(\sticky_gen.firstOne_B [2]), 
         .D(\sticky_gen.firstOne_A [2]), .Z(n39740)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i28147_4_lut.init = 16'h8228;
    LUT4 i28151_4_lut (.A(n39740), .B(n70696), .C(\sticky_gen.firstOne_B [3]), 
         .D(\sticky_gen.firstOne_A [3]), .Z(n39744)) /* synthesis lut_function=(A+(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i28151_4_lut.init = 16'hebbe;
    LUT4 i2_4_lut_adj_882 (.A(n4_adj_485), .B(n39744), .C(n8), .D(n62771), 
         .Z(n63126)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B+(C+!(D)))) */ ;
    defparam i2_4_lut_adj_882.init = 16'hd4fd;
    LUT4 i2_4_lut_adj_883 (.A(\prod[21] ), .B(n63126), .C(\prod[47] ), 
         .D(\prod[22] ), .Z(n63205)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i2_4_lut_adj_883.init = 16'hfbbb;
    LUT4 i1_4_lut_adj_884 (.A(\prod[23] ), .B(\prod[22] ), .C(\prod[24] ), 
         .D(\prod[47] ), .Z(n64329)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_884.init = 16'ha088;
    LUT4 mux_122_i18_3_lut (.A(\prod[37] ), .B(\prod[38] ), .C(\prod[47] ), 
         .Z(frac_norm[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i18_3_lut.init = 16'hcaca;
    LUT4 mux_122_i20_3_lut (.A(\prod[39] ), .B(\prod[40] ), .C(\prod[47] ), 
         .Z(frac_norm[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i20_3_lut.init = 16'hcaca;
    LUT4 mux_122_i19_3_lut (.A(\prod[38] ), .B(\prod[39] ), .C(\prod[47] ), 
         .Z(frac_norm[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i19_3_lut.init = 16'hcaca;
    LUT4 mux_122_i22_3_lut (.A(\prod[41] ), .B(\prod[42] ), .C(\prod[47] ), 
         .Z(frac_norm[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i22_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_885 (.A(\B_int[5] ), .B(\B_int[4] ), .Z(n23)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_885.init = 16'heeee;
    LUT4 mux_122_i24_3_lut (.A(\prod[43] ), .B(\prod[44] ), .C(\prod[47] ), 
         .Z(frac_norm[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i24_3_lut.init = 16'hcaca;
    LUT4 mux_122_i23_3_lut (.A(\prod[42] ), .B(\prod[43] ), .C(\prod[47] ), 
         .Z(frac_norm[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i23_3_lut.init = 16'hcaca;
    LUT4 i55133_4_lut (.A(\B_int[8] ), .B(\B_int[15] ), .C(n70839), .D(\B_int[14] ), 
         .Z(n67053)) /* synthesis lut_function=(A+!(B (C)+!B (C+!(D)))) */ ;
    defparam i55133_4_lut.init = 16'hafae;
    LUT4 mux_122_i26_3_lut (.A(\prod[45] ), .B(\prod[46] ), .C(\prod[47] ), 
         .Z(frac_norm[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i26_3_lut.init = 16'hcaca;
    LUT4 mux_122_i25_3_lut (.A(\prod[44] ), .B(\prod[45] ), .C(\prod[47] ), 
         .Z(frac_norm[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_122_i25_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_886 (.A(\B_int[0] ), .B(\B_int[1] ), .C(n12_adj_487), 
         .Z(n346[0])) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i1_3_lut_adj_886.init = 16'h5454;
    LUT4 i1_3_lut_adj_887 (.A(\B_int[14] ), .B(\B_int[15] ), .C(\B_int[16] ), 
         .Z(n16)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;
    defparam i1_3_lut_adj_887.init = 16'h4545;
    LUT4 i55134_4_lut (.A(\B_int[8] ), .B(\B_int[12] ), .C(\B_int[13] ), 
         .D(n16), .Z(n67051)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;
    defparam i55134_4_lut.init = 16'hbbba;
    
endmodule
//
// Verilog Description of module \fp_exp_clk(8,23) 
//

module \fp_exp_clk(8,23)  (clock, fR1_e3, GND_net, ufl1_e3, \fR1_e3[22] , 
            \fR1_e3[21] , \fR1_e3[20] , \fR1_e3[19] , \fR1_e3[18] , 
            \fR1_e3[17] , \fR1_e3[16] , \fR1_e3[15] , \fR1_e3[14] , 
            \fR1_e3[13] , \fR1_e3[12] , \fR1_e3[11] , \fR1_e3[10] , 
            \fR1_e3[9] , \fR1_e3[8] , \fR1_e3[7] , \fR1_e3[6] , \fR1_e3[5] , 
            \fR1_e3[4] , \fR1_e3[3] , \fR1_e3[2] , \fR1_e3[1] , \eR_e3[7] , 
            \eR_e3[5] , \eR_e3[6] , \eR_e3[3] , \eR_e3[4] , \eR_e3[1] , 
            \eR_e3[2] , \eR_e3[0] , \mXs_0[24] , \exp_a[0] , \exp_a[1] , 
            \exp_a[2] , \exp_a[3] , \exp_a[4] , \exp_a[5] , \exp_a[6] , 
            \exp_a[7] , \exp_a[8] , \exp_a[9] , \exp_a[10] , \exp_a[11] , 
            \exp_a[12] , \exp_a[13] , \exp_a[14] , \exp_a[15] , \exp_a[16] , 
            \exp_a[17] , \exp_a[18] , \exp_a[19] , \exp_a[20] , \exp_a[21] , 
            \exp_a[22] , \exp_a[30] , \exp_a[28] , \exp_a[29] , \exp_a[26] , 
            \exp_a[27] , \exp_a[24] , \exp_a[25] , \exp_a[23] , VCC_net, 
            \buf_x[89] , \buf_x[87] , \buf_x[88] , \buf_x[85] , \buf_x[86] , 
            \buf_x[83] , \buf_x[84] , \buf_r[89] , \buf_r[87] , \buf_r[88] , 
            \buf_r[85] , \buf_r[86] , \buf_r[83] , \buf_r[84] , \exp_a[32] );
    input clock;
    output [23:0]fR1_e3;
    input GND_net;
    output ufl1_e3;
    output \fR1_e3[22] ;
    output \fR1_e3[21] ;
    output \fR1_e3[20] ;
    output \fR1_e3[19] ;
    output \fR1_e3[18] ;
    output \fR1_e3[17] ;
    output \fR1_e3[16] ;
    output \fR1_e3[15] ;
    output \fR1_e3[14] ;
    output \fR1_e3[13] ;
    output \fR1_e3[12] ;
    output \fR1_e3[11] ;
    output \fR1_e3[10] ;
    output \fR1_e3[9] ;
    output \fR1_e3[8] ;
    output \fR1_e3[7] ;
    output \fR1_e3[6] ;
    output \fR1_e3[5] ;
    output \fR1_e3[4] ;
    output \fR1_e3[3] ;
    output \fR1_e3[2] ;
    output \fR1_e3[1] ;
    output \eR_e3[7] ;
    output \eR_e3[5] ;
    output \eR_e3[6] ;
    output \eR_e3[3] ;
    output \eR_e3[4] ;
    output \eR_e3[1] ;
    output \eR_e3[2] ;
    output \eR_e3[0] ;
    input \mXs_0[24] ;
    input \exp_a[0] ;
    input \exp_a[1] ;
    input \exp_a[2] ;
    input \exp_a[3] ;
    input \exp_a[4] ;
    input \exp_a[5] ;
    input \exp_a[6] ;
    input \exp_a[7] ;
    input \exp_a[8] ;
    input \exp_a[9] ;
    input \exp_a[10] ;
    input \exp_a[11] ;
    input \exp_a[12] ;
    input \exp_a[13] ;
    input \exp_a[14] ;
    input \exp_a[15] ;
    input \exp_a[16] ;
    input \exp_a[17] ;
    input \exp_a[18] ;
    input \exp_a[19] ;
    input \exp_a[20] ;
    input \exp_a[21] ;
    input \exp_a[22] ;
    input \exp_a[30] ;
    input \exp_a[28] ;
    input \exp_a[29] ;
    input \exp_a[26] ;
    input \exp_a[27] ;
    input \exp_a[24] ;
    input \exp_a[25] ;
    input \exp_a[23] ;
    input VCC_net;
    output \buf_x[89] ;
    output \buf_x[87] ;
    output \buf_x[88] ;
    output \buf_x[85] ;
    output \buf_x[86] ;
    output \buf_x[83] ;
    output \buf_x[84] ;
    input \buf_r[89] ;
    input \buf_r[87] ;
    input \buf_r[88] ;
    input \buf_r[85] ;
    input \buf_r[86] ;
    input \buf_r[83] ;
    input \buf_r[84] ;
    input \exp_a[32] ;
    
    wire ufl0_a1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(830[10:17])
    wire [0:0]nX_d;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(829[10:17])
    wire [43:0]nKLog2_c1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(793[10:19])
    wire [43:0]nKLog2_c0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(792[10:19])
    wire [20:0]nZ2_e1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(809[10:16])
    wire [49:0]nZ1_e0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(807[10:16])
    wire [27:0]nZ_e2;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(811[10:15])
    wire [27:0]nZ_e1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(810[10:15])
    wire [24:0]fR0_e2;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(818[10:16])
    wire [24:0]fR0_e1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(817[10:16])
    wire [27:0]nZ_e3;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(812[10:15])
    wire [23:0]fR1_e2;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(819[10:16])
    wire [33:0]fpX_e3;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(777[10:16])
    wire [509:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    wire [13:0]r_1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(7717[10:13])
    wire [13:0]r_0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(7709[10:13])
    wire [12:0]nEY2_d1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(803[10:17])
    wire [35:0]nY_d1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(796[10:15])
    wire [21:0]nZ0_d1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(805[10:16])
    wire [23:0]fR1_e3_c;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(820[10:16])
    wire [27:0]nEY1_e1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(801[10:17])
    wire [21:0]nK0_b0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(785[10:16])
    wire [8:0]nK_b0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(786[10:15])
    wire [35:0]nY_c1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(795[10:15])
    wire [7:0]nY1_c1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(797[10:16])
    wire [8:0]nK_e3;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(788[10:15])
    wire [11:0]eX_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(533[10:14])
    wire [35:0]nX_a0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(779[10:15])
    wire [615:0]buf_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(544[10:15])
    wire [27:0]nEY1_d2;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(800[10:17])
    wire [21:0]nZ0_d2;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(806[10:16])
    wire [1195:0]buf_x_adj_466;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [1195:0]buf_r;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(337[10:15])
    wire [35:0]nX_a1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(780[10:15])
    wire [482:0]buf_x_adj_467;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [107:0]buf_adj_468;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    wire [27:0]nEY1_c1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(799[10:17])
    wire [35:0]nX_c1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(781[10:15])
    wire [13:0]n15445;
    
    wire n70868, n65483, n62529, n14726, n62528, n62527, n62526, 
        n62525, n62524, n62523, n62522, n62521, n62520, n62519, 
        n62518, n992;
    wire [13:0]n15461;
    
    wire n17466, n62, n61502, n61501, n61500, n61499, n61664, 
        n61663, n61662, n61661, n61660, n61659, n61658, n61657, 
        n61656, n61655, n61654, n61653, n61652, n61650, n61649, 
        n61648, n61647, n61646, n61645, n61644, n61643, n61642, 
        n61641, n61639, n61638, n61637, n61636, n23965, n23964, 
        n23963, n23962, n23961, n23960, n23959, n23958, n23957, 
        n23956, n62787;
    
    FD1S3AX ufl0_a1_46 (.D(nX_d[0]), .CK(clock), .Q(ufl0_a1));
    defparam ufl0_a1_46.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i1 (.D(nKLog2_c0[7]), .CK(clock), .Q(nKLog2_c1[7]));
    defparam nKLog2_c1_i1.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i0 (.D(nZ1_e0[29]), .CK(clock), .Q(nZ2_e1[0]));
    defparam nZ2_e1_i0.GSR = "DISABLED";
    FD1S3AX nZ_e2_i1 (.D(nZ_e1[27]), .CK(clock), .Q(nZ_e2[27]));
    defparam nZ_e2_i1.GSR = "DISABLED";
    FD1S3AX fR0_e2_i0 (.D(fR0_e1[0]), .CK(clock), .Q(fR0_e2[0]));
    defparam fR0_e2_i0.GSR = "DISABLED";
    FD1S3AX nZ_e3_i1 (.D(nZ_e2[27]), .CK(clock), .Q(nZ_e3[27]));
    defparam nZ_e3_i1.GSR = "DISABLED";
    FD1S3AX fR1_e3_i0 (.D(fR1_e2[0]), .CK(clock), .Q(fR1_e3[0]));
    defparam fR1_e3_i0.GSR = "DISABLED";
    FD1S3AX buf_508__481 (.D(\buf [474]), .CK(clock), .Q(fpX_e3[32]));
    defparam buf_508__481.GSR = "DISABLED";
    FD1S3IX nEY2_d1_ret0_i12 (.D(n65483), .CK(clock), .CD(n70868), .Q(n15445[11]));
    defparam nEY2_d1_ret0_i12.GSR = "DISABLED";
    CCU2D add_4625_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62529), 
          .S0(n14726));
    defparam add_4625_cout.INIT0 = 16'h0000;
    defparam add_4625_cout.INIT1 = 16'h0000;
    defparam add_4625_cout.INJECT1_0 = "NO";
    defparam add_4625_cout.INJECT1_1 = "NO";
    CCU2D add_4625_23 (.A0(fR0_e2[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62528), .COUT(n62529), .S0(fR1_e2[21]), .S1(fR1_e2[22]));
    defparam add_4625_23.INIT0 = 16'h5aaa;
    defparam add_4625_23.INIT1 = 16'h5aaa;
    defparam add_4625_23.INJECT1_0 = "NO";
    defparam add_4625_23.INJECT1_1 = "NO";
    CCU2D add_4625_21 (.A0(fR0_e2[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62527), .COUT(n62528), .S0(fR1_e2[19]), .S1(fR1_e2[20]));
    defparam add_4625_21.INIT0 = 16'h5aaa;
    defparam add_4625_21.INIT1 = 16'h5aaa;
    defparam add_4625_21.INJECT1_0 = "NO";
    defparam add_4625_21.INJECT1_1 = "NO";
    CCU2D add_4625_19 (.A0(fR0_e2[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62526), .COUT(n62527), .S0(fR1_e2[17]), .S1(fR1_e2[18]));
    defparam add_4625_19.INIT0 = 16'h5aaa;
    defparam add_4625_19.INIT1 = 16'h5aaa;
    defparam add_4625_19.INJECT1_0 = "NO";
    defparam add_4625_19.INJECT1_1 = "NO";
    CCU2D add_4625_17 (.A0(fR0_e2[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62525), .COUT(n62526), .S0(fR1_e2[15]), .S1(fR1_e2[16]));
    defparam add_4625_17.INIT0 = 16'h5aaa;
    defparam add_4625_17.INIT1 = 16'h5aaa;
    defparam add_4625_17.INJECT1_0 = "NO";
    defparam add_4625_17.INJECT1_1 = "NO";
    CCU2D add_4625_15 (.A0(fR0_e2[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62524), .COUT(n62525), .S0(fR1_e2[13]), .S1(fR1_e2[14]));
    defparam add_4625_15.INIT0 = 16'h5aaa;
    defparam add_4625_15.INIT1 = 16'h5aaa;
    defparam add_4625_15.INJECT1_0 = "NO";
    defparam add_4625_15.INJECT1_1 = "NO";
    CCU2D add_4625_13 (.A0(fR0_e2[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62523), .COUT(n62524), .S0(fR1_e2[11]), .S1(fR1_e2[12]));
    defparam add_4625_13.INIT0 = 16'h5aaa;
    defparam add_4625_13.INIT1 = 16'h5aaa;
    defparam add_4625_13.INJECT1_0 = "NO";
    defparam add_4625_13.INJECT1_1 = "NO";
    CCU2D add_4625_11 (.A0(fR0_e2[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62522), .COUT(n62523), .S0(fR1_e2[9]), .S1(fR1_e2[10]));
    defparam add_4625_11.INIT0 = 16'h5aaa;
    defparam add_4625_11.INIT1 = 16'h5aaa;
    defparam add_4625_11.INJECT1_0 = "NO";
    defparam add_4625_11.INJECT1_1 = "NO";
    CCU2D add_4625_9 (.A0(fR0_e2[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62521), .COUT(n62522), .S0(fR1_e2[7]), .S1(fR1_e2[8]));
    defparam add_4625_9.INIT0 = 16'h5aaa;
    defparam add_4625_9.INIT1 = 16'h5aaa;
    defparam add_4625_9.INJECT1_0 = "NO";
    defparam add_4625_9.INJECT1_1 = "NO";
    CCU2D add_4625_7 (.A0(fR0_e2[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62520), .COUT(n62521), .S0(fR1_e2[5]), .S1(fR1_e2[6]));
    defparam add_4625_7.INIT0 = 16'h5aaa;
    defparam add_4625_7.INIT1 = 16'h5aaa;
    defparam add_4625_7.INJECT1_0 = "NO";
    defparam add_4625_7.INJECT1_1 = "NO";
    CCU2D add_4625_5 (.A0(fR0_e2[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62519), .COUT(n62520), .S0(fR1_e2[3]), .S1(fR1_e2[4]));
    defparam add_4625_5.INIT0 = 16'h5aaa;
    defparam add_4625_5.INIT1 = 16'h5aaa;
    defparam add_4625_5.INJECT1_0 = "NO";
    defparam add_4625_5.INJECT1_1 = "NO";
    CCU2D add_4625_3 (.A0(fR0_e2[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62518), .COUT(n62519), .S0(fR1_e2[1]), .S1(fR1_e2[2]));
    defparam add_4625_3.INIT0 = 16'h5aaa;
    defparam add_4625_3.INIT1 = 16'h5aaa;
    defparam add_4625_3.INJECT1_0 = "NO";
    defparam add_4625_3.INJECT1_1 = "NO";
    CCU2D add_4625_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(fR0_e2[1]), .B1(n992), .C1(fR0_e2[2]), .D1(GND_net), .COUT(n62518), 
          .S1(fR1_e2[0]));
    defparam add_4625_1.INIT0 = 16'hF000;
    defparam add_4625_1.INIT1 = 16'h7878;
    defparam add_4625_1.INJECT1_0 = "NO";
    defparam add_4625_1.INJECT1_1 = "NO";
    FD1S3AX nEY2_d1_ret1_i1 (.D(r_1[0]), .CK(clock), .Q(n15461[0]));
    defparam nEY2_d1_ret1_i1.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i1 (.D(r_0[0]), .CK(clock), .Q(n15445[0]));
    defparam nEY2_d1_ret0_i1.GSR = "DISABLED";
    LUT4 i49844_2_lut (.A(nEY2_d1[1]), .B(nY_d1[0]), .Z(nZ0_d1[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49844_2_lut.init = 16'h6666;
    LUT4 i27808_2_lut (.A(ufl0_a1), .B(fpX_e3[32]), .Z(ufl1_e3)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i27808_2_lut.init = 16'hbbbb;
    FD1S3AX fR1_e3_i23 (.D(n14726), .CK(clock), .Q(fR1_e3_c[23]));
    defparam fR1_e3_i23.GSR = "DISABLED";
    FD1S3AX fR1_e3_i22 (.D(fR1_e2[22]), .CK(clock), .Q(\fR1_e3[22] ));
    defparam fR1_e3_i22.GSR = "DISABLED";
    FD1S3AX fR1_e3_i21 (.D(fR1_e2[21]), .CK(clock), .Q(\fR1_e3[21] ));
    defparam fR1_e3_i21.GSR = "DISABLED";
    FD1S3AX fR1_e3_i20 (.D(fR1_e2[20]), .CK(clock), .Q(\fR1_e3[20] ));
    defparam fR1_e3_i20.GSR = "DISABLED";
    FD1S3AX fR1_e3_i19 (.D(fR1_e2[19]), .CK(clock), .Q(\fR1_e3[19] ));
    defparam fR1_e3_i19.GSR = "DISABLED";
    FD1S3AX fR1_e3_i18 (.D(fR1_e2[18]), .CK(clock), .Q(\fR1_e3[18] ));
    defparam fR1_e3_i18.GSR = "DISABLED";
    FD1S3AX fR1_e3_i17 (.D(fR1_e2[17]), .CK(clock), .Q(\fR1_e3[17] ));
    defparam fR1_e3_i17.GSR = "DISABLED";
    FD1S3AX fR1_e3_i16 (.D(fR1_e2[16]), .CK(clock), .Q(\fR1_e3[16] ));
    defparam fR1_e3_i16.GSR = "DISABLED";
    FD1S3AX fR1_e3_i15 (.D(fR1_e2[15]), .CK(clock), .Q(\fR1_e3[15] ));
    defparam fR1_e3_i15.GSR = "DISABLED";
    FD1S3AX fR1_e3_i14 (.D(fR1_e2[14]), .CK(clock), .Q(\fR1_e3[14] ));
    defparam fR1_e3_i14.GSR = "DISABLED";
    FD1S3AX fR1_e3_i13 (.D(fR1_e2[13]), .CK(clock), .Q(\fR1_e3[13] ));
    defparam fR1_e3_i13.GSR = "DISABLED";
    FD1S3AX fR1_e3_i12 (.D(fR1_e2[12]), .CK(clock), .Q(\fR1_e3[12] ));
    defparam fR1_e3_i12.GSR = "DISABLED";
    FD1S3AX fR1_e3_i11 (.D(fR1_e2[11]), .CK(clock), .Q(\fR1_e3[11] ));
    defparam fR1_e3_i11.GSR = "DISABLED";
    FD1S3AX fR1_e3_i10 (.D(fR1_e2[10]), .CK(clock), .Q(\fR1_e3[10] ));
    defparam fR1_e3_i10.GSR = "DISABLED";
    FD1S3AX fR1_e3_i9 (.D(fR1_e2[9]), .CK(clock), .Q(\fR1_e3[9] ));
    defparam fR1_e3_i9.GSR = "DISABLED";
    FD1S3AX fR1_e3_i8 (.D(fR1_e2[8]), .CK(clock), .Q(\fR1_e3[8] ));
    defparam fR1_e3_i8.GSR = "DISABLED";
    FD1S3AX fR1_e3_i7 (.D(fR1_e2[7]), .CK(clock), .Q(\fR1_e3[7] ));
    defparam fR1_e3_i7.GSR = "DISABLED";
    FD1S3AX fR1_e3_i6 (.D(fR1_e2[6]), .CK(clock), .Q(\fR1_e3[6] ));
    defparam fR1_e3_i6.GSR = "DISABLED";
    FD1S3AX fR1_e3_i5 (.D(fR1_e2[5]), .CK(clock), .Q(\fR1_e3[5] ));
    defparam fR1_e3_i5.GSR = "DISABLED";
    FD1S3AX fR1_e3_i4 (.D(fR1_e2[4]), .CK(clock), .Q(\fR1_e3[4] ));
    defparam fR1_e3_i4.GSR = "DISABLED";
    FD1S3AX fR1_e3_i3 (.D(fR1_e2[3]), .CK(clock), .Q(\fR1_e3[3] ));
    defparam fR1_e3_i3.GSR = "DISABLED";
    FD1S3AX fR1_e3_i2 (.D(fR1_e2[2]), .CK(clock), .Q(\fR1_e3[2] ));
    defparam fR1_e3_i2.GSR = "DISABLED";
    FD1S3AX fR1_e3_i1 (.D(fR1_e2[1]), .CK(clock), .Q(\fR1_e3[1] ));
    defparam fR1_e3_i1.GSR = "DISABLED";
    FD1S3AX fR0_e2_i24 (.D(fR0_e1[24]), .CK(clock), .Q(fR0_e2[24]));
    defparam fR0_e2_i24.GSR = "DISABLED";
    FD1S3AX fR0_e2_i23 (.D(fR0_e1[23]), .CK(clock), .Q(fR0_e2[23]));
    defparam fR0_e2_i23.GSR = "DISABLED";
    FD1S3AX fR0_e2_i22 (.D(fR0_e1[22]), .CK(clock), .Q(fR0_e2[22]));
    defparam fR0_e2_i22.GSR = "DISABLED";
    FD1S3AX fR0_e2_i21 (.D(fR0_e1[21]), .CK(clock), .Q(fR0_e2[21]));
    defparam fR0_e2_i21.GSR = "DISABLED";
    FD1S3AX fR0_e2_i20 (.D(fR0_e1[20]), .CK(clock), .Q(fR0_e2[20]));
    defparam fR0_e2_i20.GSR = "DISABLED";
    FD1S3AX fR0_e2_i19 (.D(fR0_e1[19]), .CK(clock), .Q(fR0_e2[19]));
    defparam fR0_e2_i19.GSR = "DISABLED";
    FD1S3AX fR0_e2_i18 (.D(fR0_e1[18]), .CK(clock), .Q(fR0_e2[18]));
    defparam fR0_e2_i18.GSR = "DISABLED";
    FD1S3AX fR0_e2_i17 (.D(fR0_e1[17]), .CK(clock), .Q(fR0_e2[17]));
    defparam fR0_e2_i17.GSR = "DISABLED";
    FD1S3AX fR0_e2_i16 (.D(fR0_e1[16]), .CK(clock), .Q(fR0_e2[16]));
    defparam fR0_e2_i16.GSR = "DISABLED";
    FD1S3AX fR0_e2_i15 (.D(fR0_e1[15]), .CK(clock), .Q(fR0_e2[15]));
    defparam fR0_e2_i15.GSR = "DISABLED";
    FD1S3AX fR0_e2_i14 (.D(fR0_e1[14]), .CK(clock), .Q(fR0_e2[14]));
    defparam fR0_e2_i14.GSR = "DISABLED";
    FD1S3AX fR0_e2_i13 (.D(fR0_e1[13]), .CK(clock), .Q(fR0_e2[13]));
    defparam fR0_e2_i13.GSR = "DISABLED";
    FD1S3AX fR0_e2_i12 (.D(fR0_e1[12]), .CK(clock), .Q(fR0_e2[12]));
    defparam fR0_e2_i12.GSR = "DISABLED";
    FD1S3AX fR0_e2_i11 (.D(fR0_e1[11]), .CK(clock), .Q(fR0_e2[11]));
    defparam fR0_e2_i11.GSR = "DISABLED";
    FD1S3AX fR0_e2_i10 (.D(fR0_e1[10]), .CK(clock), .Q(fR0_e2[10]));
    defparam fR0_e2_i10.GSR = "DISABLED";
    FD1S3AX fR0_e2_i9 (.D(fR0_e1[9]), .CK(clock), .Q(fR0_e2[9]));
    defparam fR0_e2_i9.GSR = "DISABLED";
    FD1S3AX fR0_e2_i8 (.D(fR0_e1[8]), .CK(clock), .Q(fR0_e2[8]));
    defparam fR0_e2_i8.GSR = "DISABLED";
    FD1S3AX fR0_e2_i7 (.D(fR0_e1[7]), .CK(clock), .Q(fR0_e2[7]));
    defparam fR0_e2_i7.GSR = "DISABLED";
    FD1S3AX fR0_e2_i6 (.D(fR0_e1[6]), .CK(clock), .Q(fR0_e2[6]));
    defparam fR0_e2_i6.GSR = "DISABLED";
    FD1S3AX fR0_e2_i5 (.D(fR0_e1[5]), .CK(clock), .Q(fR0_e2[5]));
    defparam fR0_e2_i5.GSR = "DISABLED";
    FD1S3AX fR0_e2_i4 (.D(fR0_e1[4]), .CK(clock), .Q(fR0_e2[4]));
    defparam fR0_e2_i4.GSR = "DISABLED";
    FD1S3AX fR0_e2_i3 (.D(fR0_e1[3]), .CK(clock), .Q(fR0_e2[3]));
    defparam fR0_e2_i3.GSR = "DISABLED";
    FD1S3AX fR0_e2_i2 (.D(fR0_e1[2]), .CK(clock), .Q(fR0_e2[2]));
    defparam fR0_e2_i2.GSR = "DISABLED";
    FD1S3AX fR0_e2_i1 (.D(fR0_e1[1]), .CK(clock), .Q(fR0_e2[1]));
    defparam fR0_e2_i1.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i20 (.D(nZ1_e0[49]), .CK(clock), .Q(nZ2_e1[20]));
    defparam nZ2_e1_i20.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i19 (.D(nZ1_e0[48]), .CK(clock), .Q(nZ2_e1[19]));
    defparam nZ2_e1_i19.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i18 (.D(nZ1_e0[47]), .CK(clock), .Q(nZ2_e1[18]));
    defparam nZ2_e1_i18.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i17 (.D(nZ1_e0[46]), .CK(clock), .Q(nZ2_e1[17]));
    defparam nZ2_e1_i17.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i16 (.D(nZ1_e0[45]), .CK(clock), .Q(nZ2_e1[16]));
    defparam nZ2_e1_i16.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i15 (.D(nZ1_e0[44]), .CK(clock), .Q(nZ2_e1[15]));
    defparam nZ2_e1_i15.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i14 (.D(nZ1_e0[43]), .CK(clock), .Q(nZ2_e1[14]));
    defparam nZ2_e1_i14.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i13 (.D(nZ1_e0[42]), .CK(clock), .Q(nZ2_e1[13]));
    defparam nZ2_e1_i13.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i12 (.D(nZ1_e0[41]), .CK(clock), .Q(nZ2_e1[12]));
    defparam nZ2_e1_i12.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i11 (.D(nZ1_e0[40]), .CK(clock), .Q(nZ2_e1[11]));
    defparam nZ2_e1_i11.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i10 (.D(nZ1_e0[39]), .CK(clock), .Q(nZ2_e1[10]));
    defparam nZ2_e1_i10.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i9 (.D(nZ1_e0[38]), .CK(clock), .Q(nZ2_e1[9]));
    defparam nZ2_e1_i9.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i8 (.D(nZ1_e0[37]), .CK(clock), .Q(nZ2_e1[8]));
    defparam nZ2_e1_i8.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i7 (.D(nZ1_e0[36]), .CK(clock), .Q(nZ2_e1[7]));
    defparam nZ2_e1_i7.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i6 (.D(nZ1_e0[35]), .CK(clock), .Q(nZ2_e1[6]));
    defparam nZ2_e1_i6.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i5 (.D(nZ1_e0[34]), .CK(clock), .Q(nZ2_e1[5]));
    defparam nZ2_e1_i5.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i4 (.D(nZ1_e0[33]), .CK(clock), .Q(nZ2_e1[4]));
    defparam nZ2_e1_i4.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i3 (.D(nZ1_e0[32]), .CK(clock), .Q(nZ2_e1[3]));
    defparam nZ2_e1_i3.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i2 (.D(nZ1_e0[31]), .CK(clock), .Q(nZ2_e1[2]));
    defparam nZ2_e1_i2.GSR = "DISABLED";
    FD1S3AX nZ2_e1_i1 (.D(nZ1_e0[30]), .CK(clock), .Q(nZ2_e1[1]));
    defparam nZ2_e1_i1.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i28 (.D(nKLog2_c0[34]), .CK(clock), .Q(nKLog2_c1[34]));
    defparam nKLog2_c1_i28.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i27 (.D(nKLog2_c0[33]), .CK(clock), .Q(nKLog2_c1[33]));
    defparam nKLog2_c1_i27.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i26 (.D(nKLog2_c0[32]), .CK(clock), .Q(nKLog2_c1[32]));
    defparam nKLog2_c1_i26.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i25 (.D(nKLog2_c0[31]), .CK(clock), .Q(nKLog2_c1[31]));
    defparam nKLog2_c1_i25.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i24 (.D(nKLog2_c0[30]), .CK(clock), .Q(nKLog2_c1[30]));
    defparam nKLog2_c1_i24.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i23 (.D(nKLog2_c0[29]), .CK(clock), .Q(nKLog2_c1[29]));
    defparam nKLog2_c1_i23.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i22 (.D(nKLog2_c0[28]), .CK(clock), .Q(nKLog2_c1[28]));
    defparam nKLog2_c1_i22.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i21 (.D(nKLog2_c0[27]), .CK(clock), .Q(nKLog2_c1[27]));
    defparam nKLog2_c1_i21.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i20 (.D(nKLog2_c0[26]), .CK(clock), .Q(nKLog2_c1[26]));
    defparam nKLog2_c1_i20.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i19 (.D(nKLog2_c0[25]), .CK(clock), .Q(nKLog2_c1[25]));
    defparam nKLog2_c1_i19.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i18 (.D(nKLog2_c0[24]), .CK(clock), .Q(nKLog2_c1[24]));
    defparam nKLog2_c1_i18.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i17 (.D(nKLog2_c0[23]), .CK(clock), .Q(nKLog2_c1[23]));
    defparam nKLog2_c1_i17.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i16 (.D(nKLog2_c0[22]), .CK(clock), .Q(nKLog2_c1[22]));
    defparam nKLog2_c1_i16.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i15 (.D(nKLog2_c0[21]), .CK(clock), .Q(nKLog2_c1[21]));
    defparam nKLog2_c1_i15.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i14 (.D(nKLog2_c0[20]), .CK(clock), .Q(nKLog2_c1[20]));
    defparam nKLog2_c1_i14.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i13 (.D(nKLog2_c0[19]), .CK(clock), .Q(nKLog2_c1[19]));
    defparam nKLog2_c1_i13.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i12 (.D(nKLog2_c0[18]), .CK(clock), .Q(nKLog2_c1[18]));
    defparam nKLog2_c1_i12.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i11 (.D(nKLog2_c0[17]), .CK(clock), .Q(nKLog2_c1[17]));
    defparam nKLog2_c1_i11.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i10 (.D(nKLog2_c0[16]), .CK(clock), .Q(nKLog2_c1[16]));
    defparam nKLog2_c1_i10.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i9 (.D(nKLog2_c0[15]), .CK(clock), .Q(nKLog2_c1[15]));
    defparam nKLog2_c1_i9.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i8 (.D(nKLog2_c0[14]), .CK(clock), .Q(nKLog2_c1[14]));
    defparam nKLog2_c1_i8.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i7 (.D(nKLog2_c0[13]), .CK(clock), .Q(nKLog2_c1[13]));
    defparam nKLog2_c1_i7.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i6 (.D(nKLog2_c0[12]), .CK(clock), .Q(nKLog2_c1[12]));
    defparam nKLog2_c1_i6.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i5 (.D(nKLog2_c0[11]), .CK(clock), .Q(nKLog2_c1[11]));
    defparam nKLog2_c1_i5.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i4 (.D(nKLog2_c0[10]), .CK(clock), .Q(nKLog2_c1[10]));
    defparam nKLog2_c1_i4.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i3 (.D(nKLog2_c0[9]), .CK(clock), .Q(nKLog2_c1[9]));
    defparam nKLog2_c1_i3.GSR = "DISABLED";
    FD1S3AX nKLog2_c1_i2 (.D(nKLog2_c0[8]), .CK(clock), .Q(nKLog2_c1[8]));
    defparam nKLog2_c1_i2.GSR = "DISABLED";
    LUT4 i6824_2_lut (.A(nZ_e1[27]), .B(nZ_e1[2]), .Z(n17466)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6824_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(nEY1_e1[0]), .B(nZ_e1[1]), .C(nZ2_e1[0]), .D(n17466), 
         .Z(fR0_e1[0])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;
    defparam i2_4_lut.init = 16'hffde;
    LUT4 i49843_2_lut (.A(nK0_b0[13]), .B(nK0_b0[12]), .Z(nK_b0[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49843_2_lut.init = 16'h6666;
    LUT4 i11_1_lut (.A(nY_c1[27]), .Z(nY1_c1[7])) /* synthesis lut_function=(!(A)) */ ;
    defparam i11_1_lut.init = 16'h5555;
    FD1S3AX nEY2_d1_ret1_i2 (.D(r_1[1]), .CK(clock), .Q(n15461[1]));
    defparam nEY2_d1_ret1_i2.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret1_i3 (.D(r_1[2]), .CK(clock), .Q(n15461[2]));
    defparam nEY2_d1_ret1_i3.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret1_i4 (.D(r_1[3]), .CK(clock), .Q(n15461[3]));
    defparam nEY2_d1_ret1_i4.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret1_i5 (.D(r_1[4]), .CK(clock), .Q(n15461[4]));
    defparam nEY2_d1_ret1_i5.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret1_i6 (.D(r_1[5]), .CK(clock), .Q(n15461[5]));
    defparam nEY2_d1_ret1_i6.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret1_i7 (.D(r_1[6]), .CK(clock), .Q(n15461[6]));
    defparam nEY2_d1_ret1_i7.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret1_i8 (.D(r_1[7]), .CK(clock), .Q(n15461[13]));
    defparam nEY2_d1_ret1_i8.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i2 (.D(r_0[1]), .CK(clock), .Q(n15445[1]));
    defparam nEY2_d1_ret0_i2.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i3 (.D(r_0[2]), .CK(clock), .Q(n15445[2]));
    defparam nEY2_d1_ret0_i3.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i4 (.D(r_0[3]), .CK(clock), .Q(n15445[3]));
    defparam nEY2_d1_ret0_i4.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i5 (.D(r_0[4]), .CK(clock), .Q(n15445[4]));
    defparam nEY2_d1_ret0_i5.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i6 (.D(r_0[5]), .CK(clock), .Q(n15445[5]));
    defparam nEY2_d1_ret0_i6.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i7 (.D(r_0[6]), .CK(clock), .Q(n15445[6]));
    defparam nEY2_d1_ret0_i7.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i8 (.D(r_0[7]), .CK(clock), .Q(n15445[7]));
    defparam nEY2_d1_ret0_i8.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i9 (.D(r_0[8]), .CK(clock), .Q(n15445[8]));
    defparam nEY2_d1_ret0_i9.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i10 (.D(r_0[9]), .CK(clock), .Q(n15445[9]));
    defparam nEY2_d1_ret0_i10.GSR = "DISABLED";
    FD1S3AX nEY2_d1_ret0_i11 (.D(r_0[10]), .CK(clock), .Q(n15445[10]));
    defparam nEY2_d1_ret0_i11.GSR = "DISABLED";
    FD1S3IX nEY2_d1_ret0_i13 (.D(n62), .CK(clock), .CD(n70868), .Q(n15445[12]));
    defparam nEY2_d1_ret0_i13.GSR = "DISABLED";
    LUT4 mux_17_i2_3_lut (.A(nZ_e1[2]), .B(nZ_e1[3]), .C(nZ_e1[27]), .Z(fR0_e1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i2_3_lut.init = 16'hcaca;
    LUT4 mux_17_i3_3_lut (.A(nZ_e1[3]), .B(nZ_e1[4]), .C(nZ_e1[27]), .Z(fR0_e1[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i3_3_lut.init = 16'hcaca;
    LUT4 mux_17_i4_3_lut (.A(nZ_e1[4]), .B(nZ_e1[5]), .C(nZ_e1[27]), .Z(fR0_e1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i4_3_lut.init = 16'hcaca;
    LUT4 mux_17_i5_3_lut (.A(nZ_e1[5]), .B(nZ_e1[6]), .C(nZ_e1[27]), .Z(fR0_e1[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i5_3_lut.init = 16'hcaca;
    LUT4 mux_17_i6_3_lut (.A(nZ_e1[6]), .B(nZ_e1[7]), .C(nZ_e1[27]), .Z(fR0_e1[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i6_3_lut.init = 16'hcaca;
    LUT4 mux_17_i7_3_lut (.A(nZ_e1[7]), .B(nZ_e1[8]), .C(nZ_e1[27]), .Z(fR0_e1[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i7_3_lut.init = 16'hcaca;
    LUT4 mux_17_i8_3_lut (.A(nZ_e1[8]), .B(nZ_e1[9]), .C(nZ_e1[27]), .Z(fR0_e1[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i8_3_lut.init = 16'hcaca;
    LUT4 mux_17_i9_3_lut (.A(nZ_e1[9]), .B(nZ_e1[10]), .C(nZ_e1[27]), 
         .Z(fR0_e1[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i9_3_lut.init = 16'hcaca;
    LUT4 mux_17_i10_3_lut (.A(nZ_e1[10]), .B(nZ_e1[11]), .C(nZ_e1[27]), 
         .Z(fR0_e1[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i10_3_lut.init = 16'hcaca;
    LUT4 mux_17_i11_3_lut (.A(nZ_e1[11]), .B(nZ_e1[12]), .C(nZ_e1[27]), 
         .Z(fR0_e1[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i11_3_lut.init = 16'hcaca;
    LUT4 mux_17_i12_3_lut (.A(nZ_e1[12]), .B(nZ_e1[13]), .C(nZ_e1[27]), 
         .Z(fR0_e1[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i12_3_lut.init = 16'hcaca;
    LUT4 mux_17_i13_3_lut (.A(nZ_e1[13]), .B(nZ_e1[14]), .C(nZ_e1[27]), 
         .Z(fR0_e1[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i13_3_lut.init = 16'hcaca;
    LUT4 mux_17_i14_3_lut (.A(nZ_e1[14]), .B(nZ_e1[15]), .C(nZ_e1[27]), 
         .Z(fR0_e1[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i14_3_lut.init = 16'hcaca;
    LUT4 mux_17_i15_3_lut (.A(nZ_e1[15]), .B(nZ_e1[16]), .C(nZ_e1[27]), 
         .Z(fR0_e1[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i15_3_lut.init = 16'hcaca;
    LUT4 mux_17_i16_3_lut (.A(nZ_e1[16]), .B(nZ_e1[17]), .C(nZ_e1[27]), 
         .Z(fR0_e1[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i16_3_lut.init = 16'hcaca;
    LUT4 mux_17_i17_3_lut (.A(nZ_e1[17]), .B(nZ_e1[18]), .C(nZ_e1[27]), 
         .Z(fR0_e1[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i17_3_lut.init = 16'hcaca;
    LUT4 mux_17_i18_3_lut (.A(nZ_e1[18]), .B(nZ_e1[19]), .C(nZ_e1[27]), 
         .Z(fR0_e1[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i18_3_lut.init = 16'hcaca;
    LUT4 mux_17_i19_3_lut (.A(nZ_e1[19]), .B(nZ_e1[20]), .C(nZ_e1[27]), 
         .Z(fR0_e1[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i19_3_lut.init = 16'hcaca;
    LUT4 mux_17_i20_3_lut (.A(nZ_e1[20]), .B(nZ_e1[21]), .C(nZ_e1[27]), 
         .Z(fR0_e1[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i20_3_lut.init = 16'hcaca;
    LUT4 mux_17_i21_3_lut (.A(nZ_e1[21]), .B(nZ_e1[22]), .C(nZ_e1[27]), 
         .Z(fR0_e1[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i21_3_lut.init = 16'hcaca;
    LUT4 mux_17_i22_3_lut (.A(nZ_e1[22]), .B(nZ_e1[23]), .C(nZ_e1[27]), 
         .Z(fR0_e1[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i22_3_lut.init = 16'hcaca;
    LUT4 mux_17_i23_3_lut (.A(nZ_e1[23]), .B(nZ_e1[24]), .C(nZ_e1[27]), 
         .Z(fR0_e1[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i23_3_lut.init = 16'hcaca;
    LUT4 mux_17_i24_3_lut (.A(nZ_e1[24]), .B(nZ_e1[25]), .C(nZ_e1[27]), 
         .Z(fR0_e1[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i24_3_lut.init = 16'hcaca;
    LUT4 mux_17_i25_3_lut (.A(nZ_e1[25]), .B(nZ_e1[26]), .C(nZ_e1[27]), 
         .Z(fR0_e1[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_17_i25_3_lut.init = 16'hcaca;
    CCU2D add_2945_9 (.A0(nK_e3[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61502), 
          .S0(\eR_e3[7] ));
    defparam add_2945_9.INIT0 = 16'h5aaa;
    defparam add_2945_9.INIT1 = 16'h0000;
    defparam add_2945_9.INJECT1_0 = "NO";
    defparam add_2945_9.INJECT1_1 = "NO";
    CCU2D add_2945_7 (.A0(nK_e3[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nK_e3[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61501), 
          .COUT(n61502), .S0(\eR_e3[5] ), .S1(\eR_e3[6] ));
    defparam add_2945_7.INIT0 = 16'h5555;
    defparam add_2945_7.INIT1 = 16'h5555;
    defparam add_2945_7.INJECT1_0 = "NO";
    defparam add_2945_7.INJECT1_1 = "NO";
    CCU2D add_2945_5 (.A0(nK_e3[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nK_e3[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61500), 
          .COUT(n61501), .S0(\eR_e3[3] ), .S1(\eR_e3[4] ));
    defparam add_2945_5.INIT0 = 16'h5555;
    defparam add_2945_5.INIT1 = 16'h5555;
    defparam add_2945_5.INJECT1_0 = "NO";
    defparam add_2945_5.INJECT1_1 = "NO";
    CCU2D add_2945_3 (.A0(nK_e3[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nK_e3[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61499), 
          .COUT(n61500), .S0(\eR_e3[1] ), .S1(\eR_e3[2] ));
    defparam add_2945_3.INIT0 = 16'h5555;
    defparam add_2945_3.INIT1 = 16'h5555;
    defparam add_2945_3.INJECT1_0 = "NO";
    defparam add_2945_3.INJECT1_1 = "NO";
    CCU2D add_2945_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nZ_e3[27]), .B1(fR1_e3_c[23]), .C1(nK_e3[0]), .D1(GND_net), 
          .COUT(n61499), .S1(\eR_e3[0] ));
    defparam add_2945_1.INIT0 = 16'hF000;
    defparam add_2945_1.INIT1 = 16'h1e1e;
    defparam add_2945_1.INJECT1_0 = "NO";
    defparam add_2945_1.INJECT1_1 = "NO";
    CCU2D add_14_28 (.A0(nEY1_e1[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61664), .S0(nZ_e1[26]), .S1(nZ_e1[27]));
    defparam add_14_28.INIT0 = 16'h5aaa;
    defparam add_14_28.INIT1 = 16'h5aaa;
    defparam add_14_28.INJECT1_0 = "NO";
    defparam add_14_28.INJECT1_1 = "NO";
    CCU2D add_14_26 (.A0(nEY1_e1[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61663), .COUT(n61664), .S0(nZ_e1[24]), .S1(nZ_e1[25]));
    defparam add_14_26.INIT0 = 16'h5aaa;
    defparam add_14_26.INIT1 = 16'h5aaa;
    defparam add_14_26.INJECT1_0 = "NO";
    defparam add_14_26.INJECT1_1 = "NO";
    CCU2D add_14_24 (.A0(nEY1_e1[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61662), .COUT(n61663), .S0(nZ_e1[22]), .S1(nZ_e1[23]));
    defparam add_14_24.INIT0 = 16'h5aaa;
    defparam add_14_24.INIT1 = 16'h5aaa;
    defparam add_14_24.INJECT1_0 = "NO";
    defparam add_14_24.INJECT1_1 = "NO";
    CCU2D add_14_22 (.A0(nEY1_e1[20]), .B0(nZ2_e1[20]), .C0(GND_net), 
          .D0(GND_net), .A1(nEY1_e1[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61661), .COUT(n61662), .S0(nZ_e1[20]), 
          .S1(nZ_e1[21]));
    defparam add_14_22.INIT0 = 16'h5666;
    defparam add_14_22.INIT1 = 16'h5aaa;
    defparam add_14_22.INJECT1_0 = "NO";
    defparam add_14_22.INJECT1_1 = "NO";
    CCU2D add_14_20 (.A0(nEY1_e1[18]), .B0(nZ2_e1[18]), .C0(GND_net), 
          .D0(GND_net), .A1(nEY1_e1[19]), .B1(nZ2_e1[19]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61660), .COUT(n61661), .S0(nZ_e1[18]), 
          .S1(nZ_e1[19]));
    defparam add_14_20.INIT0 = 16'h5666;
    defparam add_14_20.INIT1 = 16'h5666;
    defparam add_14_20.INJECT1_0 = "NO";
    defparam add_14_20.INJECT1_1 = "NO";
    CCU2D add_14_18 (.A0(nEY1_e1[16]), .B0(nZ2_e1[16]), .C0(GND_net), 
          .D0(GND_net), .A1(nEY1_e1[17]), .B1(nZ2_e1[17]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61659), .COUT(n61660), .S0(nZ_e1[16]), 
          .S1(nZ_e1[17]));
    defparam add_14_18.INIT0 = 16'h5666;
    defparam add_14_18.INIT1 = 16'h5666;
    defparam add_14_18.INJECT1_0 = "NO";
    defparam add_14_18.INJECT1_1 = "NO";
    CCU2D add_14_16 (.A0(nEY1_e1[14]), .B0(nZ2_e1[14]), .C0(GND_net), 
          .D0(GND_net), .A1(nEY1_e1[15]), .B1(nZ2_e1[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61658), .COUT(n61659), .S0(nZ_e1[14]), 
          .S1(nZ_e1[15]));
    defparam add_14_16.INIT0 = 16'h5666;
    defparam add_14_16.INIT1 = 16'h5666;
    defparam add_14_16.INJECT1_0 = "NO";
    defparam add_14_16.INJECT1_1 = "NO";
    CCU2D add_14_14 (.A0(nEY1_e1[12]), .B0(nZ2_e1[12]), .C0(GND_net), 
          .D0(GND_net), .A1(nEY1_e1[13]), .B1(nZ2_e1[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61657), .COUT(n61658), .S0(nZ_e1[12]), 
          .S1(nZ_e1[13]));
    defparam add_14_14.INIT0 = 16'h5666;
    defparam add_14_14.INIT1 = 16'h5666;
    defparam add_14_14.INJECT1_0 = "NO";
    defparam add_14_14.INJECT1_1 = "NO";
    CCU2D add_14_12 (.A0(nEY1_e1[10]), .B0(nZ2_e1[10]), .C0(GND_net), 
          .D0(GND_net), .A1(nEY1_e1[11]), .B1(nZ2_e1[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61656), .COUT(n61657), .S0(nZ_e1[10]), 
          .S1(nZ_e1[11]));
    defparam add_14_12.INIT0 = 16'h5666;
    defparam add_14_12.INIT1 = 16'h5666;
    defparam add_14_12.INJECT1_0 = "NO";
    defparam add_14_12.INJECT1_1 = "NO";
    CCU2D add_14_10 (.A0(nEY1_e1[8]), .B0(nZ2_e1[8]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[9]), .B1(nZ2_e1[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61655), .COUT(n61656), .S0(nZ_e1[8]), .S1(nZ_e1[9]));
    defparam add_14_10.INIT0 = 16'h5666;
    defparam add_14_10.INIT1 = 16'h5666;
    defparam add_14_10.INJECT1_0 = "NO";
    defparam add_14_10.INJECT1_1 = "NO";
    CCU2D add_14_8 (.A0(nEY1_e1[6]), .B0(nZ2_e1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[7]), .B1(nZ2_e1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61654), .COUT(n61655), .S0(nZ_e1[6]), .S1(nZ_e1[7]));
    defparam add_14_8.INIT0 = 16'h5666;
    defparam add_14_8.INIT1 = 16'h5666;
    defparam add_14_8.INJECT1_0 = "NO";
    defparam add_14_8.INJECT1_1 = "NO";
    CCU2D add_14_6 (.A0(nEY1_e1[4]), .B0(nZ2_e1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[5]), .B1(nZ2_e1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61653), .COUT(n61654), .S0(nZ_e1[4]), .S1(nZ_e1[5]));
    defparam add_14_6.INIT0 = 16'h5666;
    defparam add_14_6.INIT1 = 16'h5666;
    defparam add_14_6.INJECT1_0 = "NO";
    defparam add_14_6.INJECT1_1 = "NO";
    CCU2D add_14_4 (.A0(nEY1_e1[2]), .B0(nZ2_e1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[3]), .B1(nZ2_e1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61652), .COUT(n61653), .S0(nZ_e1[2]), .S1(nZ_e1[3]));
    defparam add_14_4.INIT0 = 16'h5666;
    defparam add_14_4.INIT1 = 16'h5666;
    defparam add_14_4.INJECT1_0 = "NO";
    defparam add_14_4.INJECT1_1 = "NO";
    CCU2D add_14_2 (.A0(nEY1_e1[0]), .B0(nZ2_e1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_e1[1]), .B1(nZ2_e1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61652), .S1(nZ_e1[1]));
    defparam add_14_2.INIT0 = 16'h7000;
    defparam add_14_2.INIT1 = 16'h5666;
    defparam add_14_2.INJECT1_0 = "NO";
    defparam add_14_2.INJECT1_1 = "NO";
    CCU2D add_12_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61650), 
          .S0(nZ0_d1[21]));
    defparam add_12_cout.INIT0 = 16'h0000;
    defparam add_12_cout.INIT1 = 16'h0000;
    defparam add_12_cout.INJECT1_0 = "NO";
    defparam add_12_cout.INJECT1_1 = "NO";
    CCU2D add_12_20 (.A0(nY_d1[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nY_d1[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61649), .COUT(n61650), .S0(nZ0_d1[19]), .S1(nZ0_d1[20]));
    defparam add_12_20.INIT0 = 16'hfaaa;
    defparam add_12_20.INIT1 = 16'hfaaa;
    defparam add_12_20.INJECT1_0 = "NO";
    defparam add_12_20.INJECT1_1 = "NO";
    CCU2D add_12_18 (.A0(nY_d1[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nY_d1[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61648), .COUT(n61649), .S0(nZ0_d1[17]), .S1(nZ0_d1[18]));
    defparam add_12_18.INIT0 = 16'hfaaa;
    defparam add_12_18.INIT1 = 16'hfaaa;
    defparam add_12_18.INJECT1_0 = "NO";
    defparam add_12_18.INJECT1_1 = "NO";
    CCU2D add_12_16 (.A0(nY_d1[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nY_d1[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61647), .COUT(n61648), .S0(nZ0_d1[15]), .S1(nZ0_d1[16]));
    defparam add_12_16.INIT0 = 16'hfaaa;
    defparam add_12_16.INIT1 = 16'hfaaa;
    defparam add_12_16.INJECT1_0 = "NO";
    defparam add_12_16.INJECT1_1 = "NO";
    CCU2D add_12_14 (.A0(nY_d1[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nY_d1[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61646), .COUT(n61647), .S0(nZ0_d1[13]), .S1(nZ0_d1[14]));
    defparam add_12_14.INIT0 = 16'hfaaa;
    defparam add_12_14.INIT1 = 16'hfaaa;
    defparam add_12_14.INJECT1_0 = "NO";
    defparam add_12_14.INJECT1_1 = "NO";
    CCU2D add_12_12 (.A0(nEY2_d1[11]), .B0(nY_d1[10]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY2_d1[12]), .B1(nY_d1[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61645), .COUT(n61646), .S0(nZ0_d1[11]), .S1(nZ0_d1[12]));
    defparam add_12_12.INIT0 = 16'h5666;
    defparam add_12_12.INIT1 = 16'h5666;
    defparam add_12_12.INJECT1_0 = "NO";
    defparam add_12_12.INJECT1_1 = "NO";
    CCU2D add_12_10 (.A0(nEY2_d1[9]), .B0(nY_d1[8]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY2_d1[10]), .B1(nY_d1[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61644), .COUT(n61645), .S0(nZ0_d1[9]), .S1(nZ0_d1[10]));
    defparam add_12_10.INIT0 = 16'h5666;
    defparam add_12_10.INIT1 = 16'h5666;
    defparam add_12_10.INJECT1_0 = "NO";
    defparam add_12_10.INJECT1_1 = "NO";
    CCU2D add_12_8 (.A0(nEY2_d1[7]), .B0(nY_d1[6]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY2_d1[8]), .B1(nY_d1[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61643), .COUT(n61644), .S0(nZ0_d1[7]), .S1(nZ0_d1[8]));
    defparam add_12_8.INIT0 = 16'h5666;
    defparam add_12_8.INIT1 = 16'h5666;
    defparam add_12_8.INJECT1_0 = "NO";
    defparam add_12_8.INJECT1_1 = "NO";
    CCU2D add_12_6 (.A0(nEY2_d1[5]), .B0(nY_d1[4]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY2_d1[6]), .B1(nY_d1[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61642), .COUT(n61643), .S0(nZ0_d1[5]), .S1(nZ0_d1[6]));
    defparam add_12_6.INIT0 = 16'h5666;
    defparam add_12_6.INIT1 = 16'h5666;
    defparam add_12_6.INJECT1_0 = "NO";
    defparam add_12_6.INJECT1_1 = "NO";
    CCU2D add_12_4 (.A0(nEY2_d1[3]), .B0(nY_d1[2]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY2_d1[4]), .B1(nY_d1[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61641), .COUT(n61642), .S0(nZ0_d1[3]), .S1(nZ0_d1[4]));
    defparam add_12_4.INIT0 = 16'h5666;
    defparam add_12_4.INIT1 = 16'h5666;
    defparam add_12_4.INJECT1_0 = "NO";
    defparam add_12_4.INJECT1_1 = "NO";
    CCU2D add_12_2 (.A0(nEY2_d1[1]), .B0(nY_d1[0]), .C0(GND_net), .D0(GND_net), 
          .A1(nEY2_d1[2]), .B1(nY_d1[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61641), .S1(nZ0_d1[2]));
    defparam add_12_2.INIT0 = 16'h7000;
    defparam add_12_2.INIT1 = 16'h5666;
    defparam add_12_2.INJECT1_0 = "NO";
    defparam add_12_2.INJECT1_1 = "NO";
    CCU2D add_6_10 (.A0(nK0_b0[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61639), 
          .S0(nK_b0[8]));
    defparam add_6_10.INIT0 = 16'h5aaa;
    defparam add_6_10.INIT1 = 16'h0000;
    defparam add_6_10.INJECT1_0 = "NO";
    defparam add_6_10.INJECT1_1 = "NO";
    CCU2D add_6_8 (.A0(nK0_b0[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nK0_b0[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61638), .COUT(n61639), .S0(nK_b0[6]), .S1(nK_b0[7]));
    defparam add_6_8.INIT0 = 16'h5aaa;
    defparam add_6_8.INIT1 = 16'h5aaa;
    defparam add_6_8.INJECT1_0 = "NO";
    defparam add_6_8.INJECT1_1 = "NO";
    CCU2D add_6_6 (.A0(nK0_b0[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nK0_b0[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61637), .COUT(n61638), .S0(nK_b0[4]), .S1(nK_b0[5]));
    defparam add_6_6.INIT0 = 16'h5aaa;
    defparam add_6_6.INIT1 = 16'h5aaa;
    defparam add_6_6.INJECT1_0 = "NO";
    defparam add_6_6.INJECT1_1 = "NO";
    CCU2D add_6_4 (.A0(nK0_b0[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nK0_b0[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61636), .COUT(n61637), .S0(nK_b0[2]), .S1(nK_b0[3]));
    defparam add_6_4.INIT0 = 16'h5aaa;
    defparam add_6_4.INIT1 = 16'h5aaa;
    defparam add_6_4.INJECT1_0 = "NO";
    defparam add_6_4.INJECT1_1 = "NO";
    CCU2D add_6_2 (.A0(nK0_b0[13]), .B0(nK0_b0[12]), .C0(GND_net), .D0(GND_net), 
          .A1(nK0_b0[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n61636), .S1(nK_b0[1]));
    defparam add_6_2.INIT0 = 16'h7000;
    defparam add_6_2.INIT1 = 16'h5aaa;
    defparam add_6_2.INJECT1_0 = "NO";
    defparam add_6_2.INJECT1_1 = "NO";
    LUT4 i21_2_lut (.A(fR0_e2[2]), .B(fR0_e2[0]), .Z(n992)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i21_2_lut.init = 16'heeee;
    \fp_exp_shift_clk(8,23)  shift (.clock(clock), .\eX_x[11] (eX_x[11]), 
            .\mXs_0[24] (\mXs_0[24] ), .\nX_a0[31] (nX_a0[31]), .\exp_a[0] (\exp_a[0] ), 
            .\exp_a[1] (\exp_a[1] ), .\exp_a[2] (\exp_a[2] ), .\exp_a[3] (\exp_a[3] ), 
            .\exp_a[4] (\exp_a[4] ), .\exp_a[5] (\exp_a[5] ), .\exp_a[6] (\exp_a[6] ), 
            .\exp_a[7] (\exp_a[7] ), .\exp_a[8] (\exp_a[8] ), .\exp_a[9] (\exp_a[9] ), 
            .\exp_a[10] (\exp_a[10] ), .\exp_a[11] (\exp_a[11] ), .\exp_a[12] (\exp_a[12] ), 
            .\exp_a[13] (\exp_a[13] ), .\exp_a[14] (\exp_a[14] ), .\exp_a[15] (\exp_a[15] ), 
            .\exp_a[16] (\exp_a[16] ), .\exp_a[17] (\exp_a[17] ), .\exp_a[18] (\exp_a[18] ), 
            .\exp_a[19] (\exp_a[19] ), .\exp_a[20] (\exp_a[20] ), .\exp_a[21] (\exp_a[21] ), 
            .\exp_a[22] (\exp_a[22] ), .\nX_a0[30] (nX_a0[30]), .\buf_x[463] (buf_x[463]), 
            .\exp_a[30] (\exp_a[30] ), .GND_net(GND_net), .\exp_a[28] (\exp_a[28] ), 
            .\exp_a[29] (\exp_a[29] ), .\exp_a[26] (\exp_a[26] ), .\exp_a[27] (\exp_a[27] ), 
            .\exp_a[24] (\exp_a[24] ), .\exp_a[25] (\exp_a[25] ), .\exp_a[23] (\exp_a[23] ), 
            .\buf_x[467] (buf_x[467]), .\buf_x[468] (buf_x[468]), .\buf_x[469] (buf_x[469]), 
            .\buf_x[470] (buf_x[470]), .\buf_x[471] (buf_x[471]), .\nX_a0[32] (nX_a0[32]), 
            .\buf_x[464] (buf_x[464]), .\nX_a0[33] (nX_a0[33]), .\buf_x[465] (buf_x[465]), 
            .\nX_a0[34] (nX_a0[34]), .\buf_x[466] (buf_x[466]), .\nX_a0[35] (nX_a0[35]), 
            .\nX_a0[24] (nX_a0[24]), .\nX_a0[23] (nX_a0[23]), .\nX_a0[22] (nX_a0[22]), 
            .\nX_a0[21] (nX_a0[21]), .\nX_a0[20] (nX_a0[20]), .\nX_a0[19] (nX_a0[19]), 
            .\nX_a0[18] (nX_a0[18]), .\nX_a0[17] (nX_a0[17]), .\nX_a0[16] (nX_a0[16]), 
            .\nX_a0[15] (nX_a0[15]), .\nX_a0[14] (nX_a0[14]), .\nX_a0[13] (nX_a0[13]), 
            .\nX_a0[12] (nX_a0[12]), .\nX_a0[11] (nX_a0[11]), .\nX_a0[10] (nX_a0[10]), 
            .\nX_a0[9] (nX_a0[9]), .\nX_a0[25] (nX_a0[25]), .\nX_a0[26] (nX_a0[26]), 
            .\nX_a0[27] (nX_a0[27]), .\nX_a0[28] (nX_a0[28]), .\nX_a0[29] (nX_a0[29]), 
            .nX_d({nX_d}));
    \mult_clk(28,22,false,false,0,2)  mult_z1 (.nEY1_d2({nEY1_d2}), .nZ0_d2({nZ0_d2}), 
            .GND_net(GND_net), .clock(clock), .n23965(n23965), .n23964(n23964), 
            .n23963(n23963), .n23962(n23962), .n23961(n23961), .n23960(n23960), 
            .n23959(n23959), .n23958(n23958), .n23957(n23957), .n23956(n23956), 
            .\nZ1_e0[48] (nZ1_e0[48]), .\nZ1_e0[49] (nZ1_e0[49]), .\nZ1_e0[46] (nZ1_e0[46]), 
            .\nZ1_e0[47] (nZ1_e0[47]), .\nZ1_e0[44] (nZ1_e0[44]), .\nZ1_e0[45] (nZ1_e0[45]), 
            .\nZ1_e0[42] (nZ1_e0[42]), .\nZ1_e0[43] (nZ1_e0[43]), .\nZ1_e0[40] (nZ1_e0[40]), 
            .\nZ1_e0[41] (nZ1_e0[41]), .\nZ1_e0[38] (nZ1_e0[38]), .\nZ1_e0[39] (nZ1_e0[39]), 
            .\nZ1_e0[36] (nZ1_e0[36]), .\nZ1_e0[37] (nZ1_e0[37]), .\nZ1_e0[34] (nZ1_e0[34]), 
            .\nZ1_e0[35] (nZ1_e0[35]), .\nZ1_e0[32] (nZ1_e0[32]), .\nZ1_e0[33] (nZ1_e0[33]), 
            .\nZ1_e0[30] (nZ1_e0[30]), .\nZ1_e0[31] (nZ1_e0[31]), .\nZ1_e0[29] (nZ1_e0[29]));
    \mult_clk(9,35,true,false,-1,2)  mult_klog2 (.\buf_x[623] (buf_x_adj_466[623]), 
            .clock(clock), .nK_b0({nK_b0}), .GND_net(GND_net), .\nKLog2_c0[34] (nKLog2_c0[34]), 
            .\nKLog2_c0[32] (nKLog2_c0[32]), .\nKLog2_c0[33] (nKLog2_c0[33]), 
            .\nKLog2_c0[30] (nKLog2_c0[30]), .\nKLog2_c0[31] (nKLog2_c0[31]), 
            .\nKLog2_c0[28] (nKLog2_c0[28]), .\nKLog2_c0[29] (nKLog2_c0[29]), 
            .\nKLog2_c0[26] (nKLog2_c0[26]), .\nKLog2_c0[27] (nKLog2_c0[27]), 
            .\nKLog2_c0[24] (nKLog2_c0[24]), .\nKLog2_c0[25] (nKLog2_c0[25]), 
            .\nKLog2_c0[22] (nKLog2_c0[22]), .\nKLog2_c0[23] (nKLog2_c0[23]), 
            .\nKLog2_c0[20] (nKLog2_c0[20]), .\nKLog2_c0[21] (nKLog2_c0[21]), 
            .\nKLog2_c0[18] (nKLog2_c0[18]), .\nKLog2_c0[19] (nKLog2_c0[19]), 
            .\nKLog2_c0[16] (nKLog2_c0[16]), .\nKLog2_c0[17] (nKLog2_c0[17]), 
            .\nKLog2_c0[14] (nKLog2_c0[14]), .\nKLog2_c0[15] (nKLog2_c0[15]), 
            .\nKLog2_c0[12] (nKLog2_c0[12]), .\nKLog2_c0[13] (nKLog2_c0[13]), 
            .\nKLog2_c0[10] (nKLog2_c0[10]), .\nKLog2_c0[11] (nKLog2_c0[11]), 
            .\nKLog2_c0[9] (nKLog2_c0[9]), .\buf_x[699] (buf_x_adj_466[699]), 
            .\buf_x[689] (buf_x_adj_466[689]), .\buf_x[737] (buf_x_adj_466[737]), 
            .\buf_x[727] (buf_x_adj_466[727]), .\buf_x[651] (buf_x_adj_466[651]), 
            .\buf_x[661] (buf_x_adj_466[661]), .\buf_x[613] (buf_x_adj_466[613]), 
            .\nKLog2_c0[7] (nKLog2_c0[7]), .\buf_r[936] (buf_r[936]), .\nKLog2_c0[8] (nKLog2_c0[8]));
    \mult_clk(12,10,true,false,0,3)  mult_k (.\nX_a1[0] (nX_a1[0]), .clock(clock), 
            .\eX_x[11] (eX_x[11]), .\buf_x[463] (buf_x[463]), .\buf_x[437] (buf_x_adj_467[437]), 
            .\buf_x[436] (buf_x_adj_467[436]), .\buf_x[435] (buf_x_adj_467[435]), 
            .\buf_x[434] (buf_x_adj_467[434]), .\nX_a0[35] (nX_a0[35]), 
            .\nX_a0[34] (nX_a0[34]), .\nX_a0[33] (nX_a0[33]), .\nX_a0[32] (nX_a0[32]), 
            .\nX_a0[31] (nX_a0[31]), .\nX_a0[30] (nX_a0[30]), .\nX_a0[29] (nX_a0[29]), 
            .\nX_a0[28] (nX_a0[28]), .\nX_a0[27] (nX_a0[27]), .\nX_a0[26] (nX_a0[26]), 
            .\nX_a0[25] (nX_a0[25]), .\nX_a0[24] (nX_a0[24]), .\nX_a1[23] (nX_a1[23]), 
            .\nX_a0[23] (nX_a0[23]), .\nX_a1[22] (nX_a1[22]), .\nX_a0[22] (nX_a0[22]), 
            .\nX_a1[21] (nX_a1[21]), .\nX_a0[21] (nX_a0[21]), .\nX_a1[20] (nX_a1[20]), 
            .\nX_a0[20] (nX_a0[20]), .\nX_a1[19] (nX_a1[19]), .\nX_a0[19] (nX_a0[19]), 
            .\nX_a1[18] (nX_a1[18]), .\nX_a0[18] (nX_a0[18]), .\nX_a1[17] (nX_a1[17]), 
            .\nX_a0[17] (nX_a0[17]), .\nX_a1[16] (nX_a1[16]), .\nX_a0[16] (nX_a0[16]), 
            .\nX_a1[15] (nX_a1[15]), .\nX_a0[15] (nX_a0[15]), .\nX_a1[14] (nX_a1[14]), 
            .\nX_a0[14] (nX_a0[14]), .\nX_a1[13] (nX_a1[13]), .\nX_a0[13] (nX_a0[13]), 
            .\nX_a1[12] (nX_a1[12]), .\nX_a0[12] (nX_a0[12]), .\nX_a1[11] (nX_a1[11]), 
            .\nX_a0[11] (nX_a0[11]), .\nX_a1[10] (nX_a1[10]), .\nX_a0[10] (nX_a0[10]), 
            .\nX_a1[9] (nX_a1[9]), .\nX_a0[9] (nX_a0[9]), .\nX_a1[8] (nX_a1[8]), 
            .\buf_x[471] (buf_x[471]), .\nX_a1[7] (nX_a1[7]), .\buf_x[470] (buf_x[470]), 
            .\nX_a1[6] (nX_a1[6]), .\buf_x[469] (buf_x[469]), .\nX_a1[5] (nX_a1[5]), 
            .\buf_x[468] (buf_x[468]), .\nX_a1[4] (nX_a1[4]), .\buf_x[467] (buf_x[467]), 
            .\nX_a1[3] (nX_a1[3]), .\buf_x[466] (buf_x[466]), .\nX_a1[2] (nX_a1[2]), 
            .\buf_x[465] (buf_x[465]), .\nX_a1[1] (nX_a1[1]), .\buf_x[464] (buf_x[464]), 
            .GND_net(GND_net), .\nK0_b0[21] (nK0_b0[21]), .\nK0_b0[19] (nK0_b0[19]), 
            .\nK0_b0[20] (nK0_b0[20]), .\nK0_b0[17] (nK0_b0[17]), .\nK0_b0[18] (nK0_b0[18]), 
            .\nK0_b0[15] (nK0_b0[15]), .\nK0_b0[16] (nK0_b0[16]), .\nK0_b0[13] (nK0_b0[13]), 
            .\nK0_b0[14] (nK0_b0[14]), .\nK0_b0[12] (nK0_b0[12]));
    \fp_exp_exp_y2_clk(23)  exp_y2 (.\buf[50] (buf_adj_468[50]), .\buf[51] (buf_adj_468[51]), 
            .\buf[52] (buf_adj_468[52]), .\buf[53] (buf_adj_468[53]), .\buf[54] (buf_adj_468[54]), 
            .\buf[55] (buf_adj_468[55]), .\r_0[6] (r_0[6]), .\r_0[7] (r_0[7]), 
            .\r_0[8] (r_0[8]), .n15447(n15445[12]), .n15462(n15461[13]), 
            .GND_net(GND_net), .nEY2_d1({nEY2_d1}), .n15449(n15445[10]), 
            .n15448(n15445[11]), .n15451(n15445[8]), .n15450(n15445[9]), 
            .n15453(n15445[6]), .n15469(n15461[6]), .n15452(n15445[7]), 
            .n15455(n15445[4]), .n15471(n15461[4]), .n15454(n15445[5]), 
            .n15470(n15461[5]), .n15457(n15445[2]), .n15473(n15461[2]), 
            .n15456(n15445[3]), .n15472(n15461[3]), .n15459(n15445[0]), 
            .n15475(n15461[0]), .n15458(n15445[1]), .n15474(n15461[1]), 
            .\nY_c1[8] (nY_c1[8]), .\nY_c1[13] (nY_c1[13]), .\r_1[7] (r_1[7]), 
            .clock(clock), .\r_1[6] (r_1[6]), .\r_1[5] (r_1[5]), .\r_1[4] (r_1[4]), 
            .\r_1[3] (r_1[3]), .\r_1[2] (r_1[2]), .\r_1[1] (r_1[1]), .\r_1[0] (r_1[0]), 
            .\nY_c1[20] (nY_c1[20]), .\nY_c1[21] (nY_c1[21]), .\nY_c1[22] (nY_c1[22]), 
            .\nY_c1[23] (nY_c1[23]), .\nY_c1[24] (nY_c1[24]), .\nY_c1[25] (nY_c1[25]), 
            .\nY_c1[26] (nY_c1[26]), .\nY1_c1[7] (nY1_c1[7]), .\nEY1_c1[9] (nEY1_c1[9]), 
            .\nEY1_c1[10] (nEY1_c1[10]), .\nEY1_c1[11] (nEY1_c1[11]), .\nEY1_c1[12] (nEY1_c1[12]), 
            .\nEY1_c1[13] (nEY1_c1[13]), .\nEY1_c1[14] (nEY1_c1[14]), .\nEY1_c1[15] (nEY1_c1[15]), 
            .\nEY1_c1[16] (nEY1_c1[16]), .\nEY1_c1[17] (nEY1_c1[17]), .\nEY1_c1[0] (nEY1_c1[0]), 
            .\nEY1_c1[1] (nEY1_c1[1]), .\nEY1_c1[2] (nEY1_c1[2]), .\nEY1_c1[3] (nEY1_c1[3]), 
            .\nEY1_c1[4] (nEY1_c1[4]), .\nEY1_c1[5] (nEY1_c1[5]), .\nEY1_c1[6] (nEY1_c1[6]), 
            .\nEY1_c1[7] (nEY1_c1[7]), .\nEY1_c1[8] (nEY1_c1[8]), .VCC_net(VCC_net), 
            .\nY_c1[10] (nY_c1[10]), .\nY_c1[12] (nY_c1[12]), .\nEY1_c1[19] (nEY1_c1[19]), 
            .\nEY1_c1[20] (nEY1_c1[20]), .\nEY1_c1[21] (nEY1_c1[21]), .\nEY1_c1[22] (nEY1_c1[22]), 
            .\nEY1_c1[23] (nEY1_c1[23]), .\nEY1_c1[24] (nEY1_c1[24]), .\nEY1_c1[18] (nEY1_c1[18]), 
            .\nY_c1[19] (nY_c1[19]), .\nY_c1[18] (nY_c1[18]), .\nY_c1[17] (nY_c1[17]), 
            .\nY_c1[16] (nY_c1[16]), .\nY_c1[15] (nY_c1[15]), .\nY_c1[14] (nY_c1[14]), 
            .\nY_c1[11] (nY_c1[11]), .\nY_c1[9] (nY_c1[9]), .\buf_x[89] (\buf_x[89] ), 
            .\buf_x[87] (\buf_x[87] ), .\buf_x[88] (\buf_x[88] ), .\buf_x[85] (\buf_x[85] ), 
            .\buf_x[86] (\buf_x[86] ), .\buf_x[83] (\buf_x[83] ), .\buf_x[84] (\buf_x[84] ), 
            .\buf_r[89] (\buf_r[89] ), .\buf_r[87] (\buf_r[87] ), .\buf_r[88] (\buf_r[88] ), 
            .\buf_r[85] (\buf_r[85] ), .\buf_r[86] (\buf_r[86] ), .\buf_r[83] (\buf_r[83] ), 
            .\buf_r[84] (\buf_r[84] ));
    \fp_exp_exp_y1(23)  exp_y1 (.\nX_c1[27] (nX_c1[27]), .\nKLog2_c1[34] (nKLog2_c1[34]), 
            .GND_net(GND_net), .\nY_c1[27] (nY_c1[27]), .\nX_c1[25] (nX_c1[25]), 
            .\nKLog2_c1[32] (nKLog2_c1[32]), .\nX_c1[26] (nX_c1[26]), .\nKLog2_c1[33] (nKLog2_c1[33]), 
            .\nY_c1[25] (nY_c1[25]), .\nY_c1[26] (nY_c1[26]), .\nX_c1[23] (nX_c1[23]), 
            .\nKLog2_c1[30] (nKLog2_c1[30]), .\nX_c1[24] (nX_c1[24]), .\nKLog2_c1[31] (nKLog2_c1[31]), 
            .\nY_c1[23] (nY_c1[23]), .\nY_c1[24] (nY_c1[24]), .\nX_c1[21] (nX_c1[21]), 
            .\nKLog2_c1[28] (nKLog2_c1[28]), .\nX_c1[22] (nX_c1[22]), .\nKLog2_c1[29] (nKLog2_c1[29]), 
            .\nY_c1[21] (nY_c1[21]), .\nY_c1[22] (nY_c1[22]), .\nX_c1[19] (nX_c1[19]), 
            .\nKLog2_c1[26] (nKLog2_c1[26]), .\nX_c1[20] (nX_c1[20]), .\nKLog2_c1[27] (nKLog2_c1[27]), 
            .\nY_c1[19] (nY_c1[19]), .\nY_c1[20] (nY_c1[20]), .\nX_c1[17] (nX_c1[17]), 
            .\nKLog2_c1[24] (nKLog2_c1[24]), .\nX_c1[18] (nX_c1[18]), .\nKLog2_c1[25] (nKLog2_c1[25]), 
            .\nY_c1[17] (nY_c1[17]), .\nY_c1[18] (nY_c1[18]), .\nX_c1[15] (nX_c1[15]), 
            .\nKLog2_c1[22] (nKLog2_c1[22]), .\nX_c1[16] (nX_c1[16]), .\nKLog2_c1[23] (nKLog2_c1[23]), 
            .\nY_c1[15] (nY_c1[15]), .\nY_c1[16] (nY_c1[16]), .\nX_c1[13] (nX_c1[13]), 
            .\nKLog2_c1[20] (nKLog2_c1[20]), .\nX_c1[14] (nX_c1[14]), .\nKLog2_c1[21] (nKLog2_c1[21]), 
            .\nY_c1[13] (nY_c1[13]), .\nY_c1[14] (nY_c1[14]), .\nX_c1[11] (nX_c1[11]), 
            .\nKLog2_c1[18] (nKLog2_c1[18]), .\nX_c1[12] (nX_c1[12]), .\nKLog2_c1[19] (nKLog2_c1[19]), 
            .\nY_c1[11] (nY_c1[11]), .\nY_c1[12] (nY_c1[12]), .\nX_c1[9] (nX_c1[9]), 
            .\nKLog2_c1[16] (nKLog2_c1[16]), .\nX_c1[10] (nX_c1[10]), .\nKLog2_c1[17] (nKLog2_c1[17]), 
            .\nY_c1[9] (nY_c1[9]), .\nY_c1[10] (nY_c1[10]), .\nX_c1[7] (nX_c1[7]), 
            .\nKLog2_c1[14] (nKLog2_c1[14]), .\nX_c1[8] (nX_c1[8]), .\nKLog2_c1[15] (nKLog2_c1[15]), 
            .\nY_c1[7] (nY_c1[7]), .\nY_c1[8] (nY_c1[8]), .\nX_c1[5] (nX_c1[5]), 
            .\nKLog2_c1[12] (nKLog2_c1[12]), .\nX_c1[6] (nX_c1[6]), .\nKLog2_c1[13] (nKLog2_c1[13]), 
            .\nY_c1[5] (nY_c1[5]), .\nY_c1[6] (nY_c1[6]), .\nX_c1[3] (nX_c1[3]), 
            .\nKLog2_c1[10] (nKLog2_c1[10]), .\nX_c1[4] (nX_c1[4]), .\nKLog2_c1[11] (nKLog2_c1[11]), 
            .\nY_c1[3] (nY_c1[3]), .\nY_c1[4] (nY_c1[4]), .\nX_c1[1] (nX_c1[1]), 
            .\nKLog2_c1[8] (nKLog2_c1[8]), .\nX_c1[2] (nX_c1[2]), .\nKLog2_c1[9] (nKLog2_c1[9]), 
            .\nY_c1[1] (nY_c1[1]), .\nY_c1[2] (nY_c1[2]), .\nX_c1[0] (nX_c1[0]), 
            .\nKLog2_c1[7] (nKLog2_c1[7]), .\nY_c1[0] (nY_c1[0]), .\nEY1_c1[25] (nEY1_c1[25]), 
            .n62787(n62787));
    \delay(22,1)  delay_nz0 (.nZ0_d2({nZ0_d2}), .clock(clock), .\nZ0_d1[20] (nZ0_d1[20]), 
            .\nZ0_d1[19] (nZ0_d1[19]), .\nZ0_d1[18] (nZ0_d1[18]), .\nZ0_d1[17] (nZ0_d1[17]), 
            .\nZ0_d1[16] (nZ0_d1[16]), .\nZ0_d1[15] (nZ0_d1[15]), .\nZ0_d1[14] (nZ0_d1[14]), 
            .\nZ0_d1[13] (nZ0_d1[13]), .\nZ0_d1[12] (nZ0_d1[12]), .\nZ0_d1[11] (nZ0_d1[11]), 
            .\nZ0_d1[10] (nZ0_d1[10]), .\nZ0_d1[9] (nZ0_d1[9]), .\nZ0_d1[8] (nZ0_d1[8]), 
            .\nZ0_d1[7] (nZ0_d1[7]), .\nZ0_d1[6] (nZ0_d1[6]), .\nZ0_d1[5] (nZ0_d1[5]), 
            .\nZ0_d1[4] (nZ0_d1[4]), .\nZ0_d1[3] (nZ0_d1[3]), .\nZ0_d1[2] (nZ0_d1[2]), 
            .\nZ0_d1[1] (nZ0_d1[1]), .\nEY2_d1[0] (nEY2_d1[0]), .\nZ0_d1[21] (nZ0_d1[21]), 
            .n23956(n23956), .n23957(n23957), .n23958(n23958), .n23959(n23959), 
            .n23960(n23960), .n23961(n23961), .n23962(n23962), .n23963(n23963), 
            .n23964(n23964), .n23965(n23965));
    \delay(36,2)  delay_ny (.\buf[55] (buf_adj_468[55]), .\buf[53] (buf_adj_468[53]), 
            .\buf[52] (buf_adj_468[52]), .\buf[51] (buf_adj_468[51]), .\buf[50] (buf_adj_468[50]), 
            .n65483(n65483), .\r_0[10] (r_0[10]), .\buf[54] (buf_adj_468[54]), 
            .\r_0[1] (r_0[1]), .\nY_d1[19] (nY_d1[19]), .clock(clock), 
            .\nY_d1[18] (nY_d1[18]), .\nY_d1[17] (nY_d1[17]), .\nY_d1[16] (nY_d1[16]), 
            .\nY_d1[15] (nY_d1[15]), .\nY_d1[14] (nY_d1[14]), .\nY_d1[13] (nY_d1[13]), 
            .\nY_d1[12] (nY_d1[12]), .\nY_d1[11] (nY_d1[11]), .\nY_d1[10] (nY_d1[10]), 
            .\nY_d1[9] (nY_d1[9]), .\nY_d1[8] (nY_d1[8]), .\nY_d1[7] (nY_d1[7]), 
            .\nY_d1[6] (nY_d1[6]), .\nY_d1[5] (nY_d1[5]), .\nY_d1[4] (nY_d1[4]), 
            .\nY_d1[3] (nY_d1[3]), .\nY_d1[2] (nY_d1[2]), .\nY_d1[1] (nY_d1[1]), 
            .\nY_d1[0] (nY_d1[0]), .\nY_c1[19] (nY_c1[19]), .\nY_c1[18] (nY_c1[18]), 
            .\nY_c1[17] (nY_c1[17]), .\nY_c1[16] (nY_c1[16]), .\nY_c1[15] (nY_c1[15]), 
            .\nY_c1[14] (nY_c1[14]), .\nY_c1[13] (nY_c1[13]), .\nY_c1[12] (nY_c1[12]), 
            .\nY_c1[11] (nY_c1[11]), .\nY_c1[10] (nY_c1[10]), .\nY_c1[9] (nY_c1[9]), 
            .\nY_c1[8] (nY_c1[8]), .\nY_c1[7] (nY_c1[7]), .\nY_c1[6] (nY_c1[6]), 
            .\nY_c1[5] (nY_c1[5]), .\nY_c1[4] (nY_c1[4]), .\nY_c1[3] (nY_c1[3]), 
            .\nY_c1[2] (nY_c1[2]), .\nY_c1[1] (nY_c1[1]), .\nY_c1[0] (nY_c1[0]), 
            .n62(n62), .\r_0[9] (r_0[9]), .\r_0[4] (r_0[4]), .\r_0[0] (r_0[0]), 
            .n70868(n70868), .\r_0[3] (r_0[3]), .\r_0[5] (r_0[5]), .\r_0[2] (r_0[2]));
    \delay(36,4)  delay_nx (.\nX_c1[27] (nX_c1[27]), .clock(clock), .\nX_c1[26] (nX_c1[26]), 
            .\nX_c1[25] (nX_c1[25]), .\nX_c1[24] (nX_c1[24]), .\nX_c1[23] (nX_c1[23]), 
            .\nX_c1[22] (nX_c1[22]), .\nX_c1[21] (nX_c1[21]), .\nX_c1[20] (nX_c1[20]), 
            .\nX_c1[19] (nX_c1[19]), .\nX_c1[18] (nX_c1[18]), .\nX_c1[17] (nX_c1[17]), 
            .\nX_c1[16] (nX_c1[16]), .\nX_c1[15] (nX_c1[15]), .\nX_c1[14] (nX_c1[14]), 
            .\nX_c1[13] (nX_c1[13]), .\nX_c1[12] (nX_c1[12]), .\nX_c1[11] (nX_c1[11]), 
            .\nX_c1[10] (nX_c1[10]), .\nX_c1[9] (nX_c1[9]), .\nX_c1[8] (nX_c1[8]), 
            .\nX_c1[7] (nX_c1[7]), .\nX_c1[6] (nX_c1[6]), .\nX_c1[5] (nX_c1[5]), 
            .\nX_c1[4] (nX_c1[4]), .\nX_c1[3] (nX_c1[3]), .\nX_c1[2] (nX_c1[2]), 
            .\nX_c1[1] (nX_c1[1]), .\nX_c1[0] (nX_c1[0]), .\buf_x[437] (buf_x_adj_467[437]), 
            .\buf_x[436] (buf_x_adj_467[436]), .\buf_x[435] (buf_x_adj_467[435]), 
            .\buf_x[434] (buf_x_adj_467[434]), .\nX_a1[23] (nX_a1[23]), 
            .\nX_a1[22] (nX_a1[22]), .\nX_a1[21] (nX_a1[21]), .\nX_a1[20] (nX_a1[20]), 
            .\nX_a1[19] (nX_a1[19]), .\nX_a1[18] (nX_a1[18]), .\nX_a1[17] (nX_a1[17]), 
            .\nX_a1[16] (nX_a1[16]), .\nX_a1[15] (nX_a1[15]), .\nX_a1[14] (nX_a1[14]), 
            .\nX_a1[13] (nX_a1[13]), .\nX_a1[12] (nX_a1[12]), .\nX_a1[11] (nX_a1[11]), 
            .\nX_a1[10] (nX_a1[10]), .\nX_a1[9] (nX_a1[9]), .\nX_a1[8] (nX_a1[8]), 
            .\nX_a1[7] (nX_a1[7]), .\nX_a1[6] (nX_a1[6]), .\nX_a1[5] (nX_a1[5]), 
            .\nX_a1[4] (nX_a1[4]), .\nX_a1[3] (nX_a1[3]), .\nX_a1[2] (nX_a1[2]), 
            .\nX_a1[1] (nX_a1[1]), .\nX_a1[0] (nX_a1[0]));
    \delay(9,10)  delay_nk (.\buf_r[936] (buf_r[936]), .clock(clock), .\buf_x[699] (buf_x_adj_466[699]), 
            .\nK_e3[7] (nK_e3[7]), .\nK_e3[6] (nK_e3[6]), .\nK_e3[5] (nK_e3[5]), 
            .\nK_e3[4] (nK_e3[4]), .\nK_e3[3] (nK_e3[3]), .\nK_e3[2] (nK_e3[2]), 
            .\nK_e3[1] (nK_e3[1]), .\nK_e3[0] (nK_e3[0]), .\buf_x[727] (buf_x_adj_466[727]), 
            .\buf_x[737] (buf_x_adj_466[737]), .\buf_x[689] (buf_x_adj_466[689]), 
            .\buf_x[651] (buf_x_adj_466[651]), .\buf_x[661] (buf_x_adj_466[661]), 
            .\buf_x[613] (buf_x_adj_466[613]), .\buf_x[623] (buf_x_adj_466[623]));
    \delay(28,3)  delay_ney1_1 (.nEY1_e1({nEY1_e1}), .clock(clock), .nEY1_d2({nEY1_d2}));
    \delay(28,3)_U25  delay_ney1_0 (.nEY1_d2({nEY1_d2}), .clock(clock), 
            .\nEY1_c1[24] (nEY1_c1[24]), .\nEY1_c1[23] (nEY1_c1[23]), .\nEY1_c1[22] (nEY1_c1[22]), 
            .\nEY1_c1[21] (nEY1_c1[21]), .\nEY1_c1[20] (nEY1_c1[20]), .\nEY1_c1[19] (nEY1_c1[19]), 
            .\nEY1_c1[18] (nEY1_c1[18]), .\nEY1_c1[17] (nEY1_c1[17]), .\nEY1_c1[16] (nEY1_c1[16]), 
            .\nEY1_c1[15] (nEY1_c1[15]), .\nEY1_c1[14] (nEY1_c1[14]), .\nEY1_c1[13] (nEY1_c1[13]), 
            .\nEY1_c1[12] (nEY1_c1[12]), .\nEY1_c1[11] (nEY1_c1[11]), .\nEY1_c1[10] (nEY1_c1[10]), 
            .\nEY1_c1[9] (nEY1_c1[9]), .\nEY1_c1[8] (nEY1_c1[8]), .\nEY1_c1[7] (nEY1_c1[7]), 
            .\nEY1_c1[6] (nEY1_c1[6]), .\nEY1_c1[5] (nEY1_c1[5]), .\nEY1_c1[4] (nEY1_c1[4]), 
            .\nEY1_c1[3] (nEY1_c1[3]), .\nEY1_c1[2] (nEY1_c1[2]), .\nEY1_c1[1] (nEY1_c1[1]), 
            .\nEY1_c1[0] (nEY1_c1[0]), .\nY1_c1[7] (nY1_c1[7]), .\nY_c1[27] (nY_c1[27]), 
            .n62787(n62787), .\nEY1_c1[25] (nEY1_c1[25]));
    \delay(34,14)  delay_fpx (.\buf[474] (\buf [474]), .clock(clock), .\exp_a[32] (\exp_a[32] ));
    
endmodule
//
// Verilog Description of module \fp_exp_shift_clk(8,23) 
//

module \fp_exp_shift_clk(8,23)  (clock, \eX_x[11] , \mXs_0[24] , \nX_a0[31] , 
            \exp_a[0] , \exp_a[1] , \exp_a[2] , \exp_a[3] , \exp_a[4] , 
            \exp_a[5] , \exp_a[6] , \exp_a[7] , \exp_a[8] , \exp_a[9] , 
            \exp_a[10] , \exp_a[11] , \exp_a[12] , \exp_a[13] , \exp_a[14] , 
            \exp_a[15] , \exp_a[16] , \exp_a[17] , \exp_a[18] , \exp_a[19] , 
            \exp_a[20] , \exp_a[21] , \exp_a[22] , \nX_a0[30] , \buf_x[463] , 
            \exp_a[30] , GND_net, \exp_a[28] , \exp_a[29] , \exp_a[26] , 
            \exp_a[27] , \exp_a[24] , \exp_a[25] , \exp_a[23] , \buf_x[467] , 
            \buf_x[468] , \buf_x[469] , \buf_x[470] , \buf_x[471] , 
            \nX_a0[32] , \buf_x[464] , \nX_a0[33] , \buf_x[465] , \nX_a0[34] , 
            \buf_x[466] , \nX_a0[35] , \nX_a0[24] , \nX_a0[23] , \nX_a0[22] , 
            \nX_a0[21] , \nX_a0[20] , \nX_a0[19] , \nX_a0[18] , \nX_a0[17] , 
            \nX_a0[16] , \nX_a0[15] , \nX_a0[14] , \nX_a0[13] , \nX_a0[12] , 
            \nX_a0[11] , \nX_a0[10] , \nX_a0[9] , \nX_a0[25] , \nX_a0[26] , 
            \nX_a0[27] , \nX_a0[28] , \nX_a0[29] , nX_d);
    input clock;
    output \eX_x[11] ;
    input \mXs_0[24] ;
    output \nX_a0[31] ;
    input \exp_a[0] ;
    input \exp_a[1] ;
    input \exp_a[2] ;
    input \exp_a[3] ;
    input \exp_a[4] ;
    input \exp_a[5] ;
    input \exp_a[6] ;
    input \exp_a[7] ;
    input \exp_a[8] ;
    input \exp_a[9] ;
    input \exp_a[10] ;
    input \exp_a[11] ;
    input \exp_a[12] ;
    input \exp_a[13] ;
    input \exp_a[14] ;
    input \exp_a[15] ;
    input \exp_a[16] ;
    input \exp_a[17] ;
    input \exp_a[18] ;
    input \exp_a[19] ;
    input \exp_a[20] ;
    input \exp_a[21] ;
    input \exp_a[22] ;
    output \nX_a0[30] ;
    output \buf_x[463] ;
    input \exp_a[30] ;
    input GND_net;
    input \exp_a[28] ;
    input \exp_a[29] ;
    input \exp_a[26] ;
    input \exp_a[27] ;
    input \exp_a[24] ;
    input \exp_a[25] ;
    input \exp_a[23] ;
    output \buf_x[467] ;
    output \buf_x[468] ;
    output \buf_x[469] ;
    output \buf_x[470] ;
    output \buf_x[471] ;
    output \nX_a0[32] ;
    output \buf_x[464] ;
    output \nX_a0[33] ;
    output \buf_x[465] ;
    output \nX_a0[34] ;
    output \buf_x[466] ;
    output \nX_a0[35] ;
    output \nX_a0[24] ;
    output \nX_a0[23] ;
    output \nX_a0[22] ;
    output \nX_a0[21] ;
    output \nX_a0[20] ;
    output \nX_a0[19] ;
    output \nX_a0[18] ;
    output \nX_a0[17] ;
    output \nX_a0[16] ;
    output \nX_a0[15] ;
    output \nX_a0[14] ;
    output \nX_a0[13] ;
    output \nX_a0[12] ;
    output \nX_a0[11] ;
    output \nX_a0[10] ;
    output \nX_a0[9] ;
    output \nX_a0[25] ;
    output \nX_a0[26] ;
    output \nX_a0[27] ;
    output \nX_a0[28] ;
    output \nX_a0[29] ;
    output [0:0]nX_d;
    
    wire [9:0]eX_0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(532[10:14])
    wire [615:0]buf_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(544[10:15])
    wire [24:0]mXs_0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(542[10:15])
    wire [87:0]buf_r;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(545[10:15])
    wire [11:0]eX_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(533[10:14])
    
    wire n41530, n70794, n70746, n40725, n70764, n14083, n69079, 
        n70807, n69010, n70806, n70881, n70882, n70878, n70879, 
        n70795, n41668, n4, n69016;
    wire [22:0]n14059;
    
    wire n70875, n70876, n69147, n61695, n61694, n61693, n61692, 
        n69021, n69008, n69004, n70944, n70945, n70941, n70942, 
        n70938, n70939, n70935, n70936, n61634, n70932, n70933, 
        n61633, n61632, n70929, n70930, n70926, n70927, n61631, 
        n61630, n61629, n70920, n70921, n61628, n70917, n70918, 
        n61627, n61626, n70914, n70915, n70911, n70912, n70908, 
        n70909, n70905, n70906, n70902, n70903, n61625, n61624, 
        n61623, n70899, n70900, n70896, n70897, n70893, n70894, 
        n70890, n70891, n70887, n70888, n70884, n70885;
    
    LUT4 i29935_2_lut_3_lut (.A(eX_0[1]), .B(eX_0[2]), .C(eX_0[3]), .Z(n41530)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i29935_2_lut_3_lut.init = 16'hfefe;
    LUT4 i29138_2_lut_rep_824 (.A(eX_0[1]), .B(eX_0[2]), .Z(n70794)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i29138_2_lut_rep_824.init = 16'heeee;
    LUT4 i133_4_lut_4_lut (.A(eX_0[3]), .B(n70746), .C(buf_x[272]), .D(mXs_0[0]), 
         .Z(buf_x[360])) /* synthesis lut_function=(!(A (B+!(D))+!A !(C))) */ ;
    defparam i133_4_lut_4_lut.init = 16'h7250;
    FD1S3AX buf_r_38__329 (.D(buf_x[390]), .CK(clock), .Q(buf_r[38]));
    defparam buf_r_38__329.GSR = "DISABLED";
    FD1S3AX buf_r_37__330 (.D(buf_x[389]), .CK(clock), .Q(buf_r[37]));
    defparam buf_r_37__330.GSR = "DISABLED";
    FD1S3AX buf_r_36__331 (.D(buf_x[388]), .CK(clock), .Q(buf_r[36]));
    defparam buf_r_36__331.GSR = "DISABLED";
    FD1S3AX buf_r_35__332 (.D(buf_x[387]), .CK(clock), .Q(buf_r[35]));
    defparam buf_r_35__332.GSR = "DISABLED";
    FD1S3AX buf_r_34__333 (.D(buf_x[386]), .CK(clock), .Q(buf_r[34]));
    defparam buf_r_34__333.GSR = "DISABLED";
    FD1S3AX buf_r_33__334 (.D(buf_x[385]), .CK(clock), .Q(buf_r[33]));
    defparam buf_r_33__334.GSR = "DISABLED";
    FD1S3AX buf_r_32__335 (.D(buf_x[384]), .CK(clock), .Q(buf_r[32]));
    defparam buf_r_32__335.GSR = "DISABLED";
    FD1S3AX buf_r_31__336 (.D(buf_x[383]), .CK(clock), .Q(buf_r[31]));
    defparam buf_r_31__336.GSR = "DISABLED";
    FD1S3AX buf_r_30__337 (.D(buf_x[382]), .CK(clock), .Q(buf_r[30]));
    defparam buf_r_30__337.GSR = "DISABLED";
    FD1S3AX buf_r_29__338 (.D(buf_x[381]), .CK(clock), .Q(buf_r[29]));
    defparam buf_r_29__338.GSR = "DISABLED";
    FD1S3AX buf_r_28__339 (.D(buf_x[380]), .CK(clock), .Q(buf_r[28]));
    defparam buf_r_28__339.GSR = "DISABLED";
    FD1S3AX buf_r_27__340 (.D(buf_x[379]), .CK(clock), .Q(buf_r[27]));
    defparam buf_r_27__340.GSR = "DISABLED";
    FD1S3AX buf_r_26__341 (.D(buf_x[378]), .CK(clock), .Q(buf_r[26]));
    defparam buf_r_26__341.GSR = "DISABLED";
    FD1S3AX buf_r_25__342 (.D(buf_x[377]), .CK(clock), .Q(buf_r[25]));
    defparam buf_r_25__342.GSR = "DISABLED";
    FD1S3AX buf_r_24__343 (.D(buf_x[376]), .CK(clock), .Q(buf_r[24]));
    defparam buf_r_24__343.GSR = "DISABLED";
    FD1S3AX buf_r_23__344 (.D(buf_x[375]), .CK(clock), .Q(buf_r[23]));
    defparam buf_r_23__344.GSR = "DISABLED";
    FD1S3AX buf_r_22__345 (.D(buf_x[374]), .CK(clock), .Q(buf_r[22]));
    defparam buf_r_22__345.GSR = "DISABLED";
    FD1S3AX buf_r_21__346 (.D(buf_x[373]), .CK(clock), .Q(buf_r[21]));
    defparam buf_r_21__346.GSR = "DISABLED";
    FD1S3AX buf_r_20__347 (.D(buf_x[372]), .CK(clock), .Q(buf_r[20]));
    defparam buf_r_20__347.GSR = "DISABLED";
    FD1S3AX buf_r_19__348 (.D(buf_x[371]), .CK(clock), .Q(buf_r[19]));
    defparam buf_r_19__348.GSR = "DISABLED";
    FD1S3AX buf_r_18__349 (.D(buf_x[370]), .CK(clock), .Q(buf_r[18]));
    defparam buf_r_18__349.GSR = "DISABLED";
    FD1S3AX buf_r_17__350 (.D(buf_x[369]), .CK(clock), .Q(buf_r[17]));
    defparam buf_r_17__350.GSR = "DISABLED";
    FD1S3AX buf_r_16__351 (.D(buf_x[368]), .CK(clock), .Q(buf_r[16]));
    defparam buf_r_16__351.GSR = "DISABLED";
    FD1S3AX buf_r_15__352 (.D(buf_x[367]), .CK(clock), .Q(buf_r[15]));
    defparam buf_r_15__352.GSR = "DISABLED";
    FD1S3AX buf_r_14__353 (.D(buf_x[366]), .CK(clock), .Q(buf_r[14]));
    defparam buf_r_14__353.GSR = "DISABLED";
    FD1S3AX buf_r_13__354 (.D(buf_x[365]), .CK(clock), .Q(buf_r[13]));
    defparam buf_r_13__354.GSR = "DISABLED";
    FD1S3AX buf_r_12__355 (.D(buf_x[364]), .CK(clock), .Q(buf_r[12]));
    defparam buf_r_12__355.GSR = "DISABLED";
    FD1S3AX buf_r_11__356 (.D(buf_x[363]), .CK(clock), .Q(buf_r[11]));
    defparam buf_r_11__356.GSR = "DISABLED";
    FD1S3AX buf_r_10__357 (.D(buf_x[362]), .CK(clock), .Q(buf_r[10]));
    defparam buf_r_10__357.GSR = "DISABLED";
    FD1S3AX buf_r_9__358 (.D(buf_x[361]), .CK(clock), .Q(buf_r[9]));
    defparam buf_r_9__358.GSR = "DISABLED";
    FD1S3AX buf_r_8__359 (.D(buf_x[360]), .CK(clock), .Q(buf_r[8]));
    defparam buf_r_8__359.GSR = "DISABLED";
    FD1S3IX buf_r_7__360 (.D(buf_x[271]), .CK(clock), .CD(eX_0[3]), .Q(buf_r[7]));
    defparam buf_r_7__360.GSR = "DISABLED";
    FD1S3IX buf_r_6__361 (.D(buf_x[270]), .CK(clock), .CD(eX_0[3]), .Q(buf_r[6]));
    defparam buf_r_6__361.GSR = "DISABLED";
    FD1S3IX buf_r_5__362 (.D(buf_x[269]), .CK(clock), .CD(eX_0[3]), .Q(buf_r[5]));
    defparam buf_r_5__362.GSR = "DISABLED";
    FD1S3IX buf_r_4__363 (.D(buf_x[268]), .CK(clock), .CD(eX_0[3]), .Q(buf_r[4]));
    defparam buf_r_4__363.GSR = "DISABLED";
    FD1S3IX buf_r_2__365 (.D(buf_x[178]), .CK(clock), .CD(n40725), .Q(buf_r[2]));
    defparam buf_r_2__365.GSR = "DISABLED";
    FD1S3AX eX_r_11__368 (.D(eX_0[5]), .CK(clock), .Q(\eX_x[11] ));
    defparam eX_r_11__368.GSR = "DISABLED";
    FD1S3AX eX_r_10__369 (.D(eX_0[4]), .CK(clock), .Q(eX_x[10]));
    defparam eX_r_10__369.GSR = "DISABLED";
    FD1S3AX buf_r_39__328 (.D(\mXs_0[24] ), .CK(clock), .Q(buf_x[615]));
    defparam buf_r_39__328.GSR = "DISABLED";
    LUT4 i29941_2_lut_rep_794_3_lut (.A(eX_0[0]), .B(eX_0[1]), .C(eX_0[2]), 
         .Z(n70764)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i29941_2_lut_rep_794_3_lut.init = 16'h8080;
    LUT4 buf_x_198__bdd_3_lut_4_lut (.A(eX_0[0]), .B(eX_0[1]), .C(n14083), 
         .D(\mXs_0[24] ), .Z(n69079)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (D)) */ ;
    defparam buf_x_198__bdd_3_lut_4_lut.init = 16'hf788;
    LUT4 i29145_2_lut_rep_837 (.A(eX_0[0]), .B(eX_0[1]), .Z(n70807)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29145_2_lut_rep_837.init = 16'h8888;
    LUT4 buf_x_285__bdd_3_lut_4_lut (.A(eX_0[1]), .B(eX_0[2]), .C(\mXs_0[24] ), 
         .D(buf_x[111]), .Z(n69010)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam buf_x_285__bdd_3_lut_4_lut.init = 16'hf870;
    LUT4 i29140_2_lut_rep_836 (.A(eX_0[1]), .B(eX_0[2]), .Z(n70806)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29140_2_lut_rep_836.init = 16'h8888;
    LUT4 i6902_3_lut_4_lut (.A(eX_0[2]), .B(eX_0[3]), .C(\mXs_0[24] ), 
         .D(buf_x[199]), .Z(buf_x[387])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam i6902_3_lut_4_lut.init = 16'hf870;
    LUT4 i6900_3_lut_4_lut (.A(eX_0[2]), .B(eX_0[3]), .C(\mXs_0[24] ), 
         .D(buf_x[200]), .Z(buf_x[388])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam i6900_3_lut_4_lut.init = 16'hf870;
    LUT4 i46_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[111]), .C(buf_x[109]), 
         .Z(buf_x[199])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i46_3_lut_3_lut.init = 16'he4e4;
    LUT4 i47_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[110]), .C(buf_x[108]), 
         .Z(buf_x[198])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i47_3_lut_3_lut.init = 16'he4e4;
    LUT4 i48_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[109]), .C(buf_x[107]), 
         .Z(buf_x[197])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i48_3_lut_3_lut.init = 16'he4e4;
    LUT4 i77_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[200]), .C(buf_x[196]), 
         .Z(buf_x[288])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i77_3_lut_3_lut.init = 16'he4e4;
    LUT4 i49_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[108]), .C(buf_x[106]), 
         .Z(buf_x[196])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i49_3_lut_3_lut.init = 16'he4e4;
    LUT4 i78_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[199]), .C(buf_x[195]), 
         .Z(buf_x[287])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i78_3_lut_3_lut.init = 16'he4e4;
    LUT4 i50_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[107]), .C(buf_x[105]), 
         .Z(buf_x[195])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i50_3_lut_3_lut.init = 16'he4e4;
    LUT4 i54640_else_3_lut (.A(buf_x[615]), .B(buf_r[36]), .C(eX_x[10]), 
         .Z(n70881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54640_else_3_lut.init = 16'hcaca;
    LUT4 i54640_then_3_lut (.A(buf_r[4]), .B(buf_r[20]), .C(eX_x[10]), 
         .Z(n70882)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54640_then_3_lut.init = 16'hacac;
    PFUMX i56082 (.BLUT(n70878), .ALUT(n70879), .C0(\eX_x[11] ), .Z(\nX_a0[31] ));
    LUT4 i79_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[198]), .C(buf_x[194]), 
         .Z(buf_x[286])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i79_3_lut_3_lut.init = 16'he4e4;
    LUT4 i51_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[106]), .C(buf_x[104]), 
         .Z(buf_x[194])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i51_3_lut_3_lut.init = 16'he4e4;
    LUT4 i80_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[197]), .C(buf_x[193]), 
         .Z(buf_x[285])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i80_3_lut_3_lut.init = 16'he4e4;
    LUT4 i52_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[105]), .C(buf_x[103]), 
         .Z(buf_x[193])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i52_3_lut_3_lut.init = 16'he4e4;
    LUT4 i81_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[196]), .C(buf_x[192]), 
         .Z(buf_x[284])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i81_3_lut_3_lut.init = 16'he4e4;
    LUT4 i53_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[104]), .C(buf_x[102]), 
         .Z(buf_x[192])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i53_3_lut_3_lut.init = 16'he4e4;
    LUT4 i82_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[195]), .C(buf_x[191]), 
         .Z(buf_x[283])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i82_3_lut_3_lut.init = 16'he4e4;
    LUT4 i54_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[103]), .C(buf_x[101]), 
         .Z(buf_x[191])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i54_3_lut_3_lut.init = 16'he4e4;
    LUT4 i115_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[290]), .C(buf_x[282]), 
         .Z(buf_x[378])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i115_3_lut_3_lut.init = 16'he4e4;
    LUT4 i83_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[194]), .C(buf_x[190]), 
         .Z(buf_x[282])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i83_3_lut_3_lut.init = 16'he4e4;
    LUT4 i55_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[102]), .C(buf_x[100]), 
         .Z(buf_x[190])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i55_3_lut_3_lut.init = 16'he4e4;
    LUT4 i116_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[289]), .C(buf_x[281]), 
         .Z(buf_x[377])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i116_3_lut_3_lut.init = 16'he4e4;
    LUT4 i84_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[193]), .C(buf_x[189]), 
         .Z(buf_x[281])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i84_3_lut_3_lut.init = 16'he4e4;
    LUT4 i56_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[101]), .C(buf_x[99]), 
         .Z(buf_x[189])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i56_3_lut_3_lut.init = 16'he4e4;
    LUT4 i117_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[288]), .C(buf_x[280]), 
         .Z(buf_x[376])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i117_3_lut_3_lut.init = 16'he4e4;
    LUT4 i85_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[192]), .C(buf_x[188]), 
         .Z(buf_x[280])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i85_3_lut_3_lut.init = 16'he4e4;
    LUT4 i57_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[100]), .C(buf_x[98]), 
         .Z(buf_x[188])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i57_3_lut_3_lut.init = 16'he4e4;
    LUT4 i118_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[287]), .C(buf_x[279]), 
         .Z(buf_x[375])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i118_3_lut_3_lut.init = 16'he4e4;
    LUT4 i86_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[191]), .C(buf_x[187]), 
         .Z(buf_x[279])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i86_3_lut_3_lut.init = 16'he4e4;
    LUT4 i58_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[99]), .C(buf_x[97]), .Z(buf_x[187])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i58_3_lut_3_lut.init = 16'he4e4;
    LUT4 i119_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[286]), .C(buf_x[278]), 
         .Z(buf_x[374])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i119_3_lut_3_lut.init = 16'he4e4;
    LUT4 i87_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[190]), .C(buf_x[186]), 
         .Z(buf_x[278])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i87_3_lut_3_lut.init = 16'he4e4;
    LUT4 i59_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[98]), .C(buf_x[96]), .Z(buf_x[186])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i59_3_lut_3_lut.init = 16'he4e4;
    LUT4 i120_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[285]), .C(buf_x[277]), 
         .Z(buf_x[373])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i120_3_lut_3_lut.init = 16'he4e4;
    LUT4 i88_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[189]), .C(buf_x[185]), 
         .Z(buf_x[277])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i88_3_lut_3_lut.init = 16'he4e4;
    LUT4 i60_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[97]), .C(buf_x[95]), .Z(buf_x[185])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i60_3_lut_3_lut.init = 16'he4e4;
    LUT4 i121_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[284]), .C(buf_x[276]), 
         .Z(buf_x[372])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i121_3_lut_3_lut.init = 16'he4e4;
    LUT4 i89_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[188]), .C(buf_x[184]), 
         .Z(buf_x[276])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i89_3_lut_3_lut.init = 16'he4e4;
    LUT4 i61_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[96]), .C(buf_x[94]), .Z(buf_x[184])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i61_3_lut_3_lut.init = 16'he4e4;
    LUT4 i122_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[283]), .C(buf_x[275]), 
         .Z(buf_x[371])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i122_3_lut_3_lut.init = 16'he4e4;
    LUT4 i90_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[187]), .C(buf_x[183]), 
         .Z(buf_x[275])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i90_3_lut_3_lut.init = 16'he4e4;
    LUT4 i62_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[95]), .C(buf_x[93]), .Z(buf_x[183])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i62_3_lut_3_lut.init = 16'he4e4;
    LUT4 i123_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[282]), .C(buf_x[274]), 
         .Z(buf_x[370])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i123_3_lut_3_lut.init = 16'he4e4;
    LUT4 i91_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[186]), .C(buf_x[182]), 
         .Z(buf_x[274])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i91_3_lut_3_lut.init = 16'he4e4;
    LUT4 i63_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[94]), .C(buf_x[92]), .Z(buf_x[182])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i63_3_lut_3_lut.init = 16'he4e4;
    LUT4 i124_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[281]), .C(buf_x[273]), 
         .Z(buf_x[369])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i124_3_lut_3_lut.init = 16'he4e4;
    LUT4 i92_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[185]), .C(buf_x[181]), 
         .Z(buf_x[273])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i92_3_lut_3_lut.init = 16'he4e4;
    LUT4 i64_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[93]), .C(buf_x[91]), .Z(buf_x[181])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i64_3_lut_3_lut.init = 16'he4e4;
    LUT4 i125_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[280]), .C(buf_x[272]), 
         .Z(buf_x[368])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i125_3_lut_3_lut.init = 16'he4e4;
    LUT4 i93_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[184]), .C(buf_x[180]), 
         .Z(buf_x[272])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i93_3_lut_3_lut.init = 16'he4e4;
    LUT4 i65_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[92]), .C(buf_x[90]), .Z(buf_x[180])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i65_3_lut_3_lut.init = 16'he4e4;
    LUT4 i126_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[279]), .C(buf_x[271]), 
         .Z(buf_x[367])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i126_3_lut_3_lut.init = 16'he4e4;
    LUT4 i94_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[183]), .C(buf_x[179]), 
         .Z(buf_x[271])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i94_3_lut_3_lut.init = 16'he4e4;
    LUT4 i66_3_lut_3_lut (.A(eX_0[1]), .B(buf_x[91]), .C(buf_x[89]), .Z(buf_x[179])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i66_3_lut_3_lut.init = 16'he4e4;
    LUT4 i127_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[278]), .C(buf_x[270]), 
         .Z(buf_x[366])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i127_3_lut_3_lut.init = 16'he4e4;
    LUT4 i95_3_lut_3_lut (.A(eX_0[2]), .B(buf_x[182]), .C(buf_x[178]), 
         .Z(buf_x[270])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i95_3_lut_3_lut.init = 16'he4e4;
    LUT4 i128_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[277]), .C(buf_x[269]), 
         .Z(buf_x[365])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i128_3_lut_3_lut.init = 16'he4e4;
    LUT4 i96_4_lut_4_lut (.A(eX_0[1]), .B(eX_0[2]), .C(buf_x[181]), .D(buf_x[89]), 
         .Z(buf_x[269])) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;
    defparam i96_4_lut_4_lut.init = 16'h7430;
    LUT4 i129_3_lut_3_lut (.A(eX_0[3]), .B(buf_x[276]), .C(buf_x[268]), 
         .Z(buf_x[364])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i129_3_lut_3_lut.init = 16'he4e4;
    LUT4 i97_4_lut_4_lut (.A(eX_0[2]), .B(n70795), .C(buf_x[180]), .D(mXs_0[0]), 
         .Z(buf_x[268])) /* synthesis lut_function=(!(A (B+!(D))+!A !(C))) */ ;
    defparam i97_4_lut_4_lut.init = 16'h7250;
    LUT4 i30068_2_lut_3_lut_4_lut (.A(eX_0[0]), .B(eX_0[1]), .C(eX_0[3]), 
         .D(eX_0[2]), .Z(n41668)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30068_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i29939_2_lut_rep_776_3_lut (.A(eX_0[0]), .B(eX_0[1]), .C(eX_0[2]), 
         .Z(n70746)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i29939_2_lut_rep_776_3_lut.init = 16'hfefe;
    LUT4 i29143_2_lut_rep_825 (.A(eX_0[0]), .B(eX_0[1]), .Z(n70795)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i29143_2_lut_rep_825.init = 16'heeee;
    LUT4 i131_4_lut_4_lut (.A(eX_0[2]), .B(eX_0[3]), .C(buf_x[274]), .D(buf_x[178]), 
         .Z(buf_x[362])) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;
    defparam i131_4_lut_4_lut.init = 16'h7430;
    LUT4 i130_4_lut_4_lut (.A(eX_0[2]), .B(eX_0[3]), .C(buf_x[275]), .D(buf_x[179]), 
         .Z(buf_x[363])) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;
    defparam i130_4_lut_4_lut.init = 16'h7430;
    LUT4 i132_4_lut_4_lut (.A(eX_0[3]), .B(n70794), .C(buf_x[273]), .D(buf_x[89]), 
         .Z(buf_x[361])) /* synthesis lut_function=(!(A (B+!(D))+!A !(C))) */ ;
    defparam i132_4_lut_4_lut.init = 16'h7250;
    LUT4 i4_1_lut (.A(n4), .Z(eX_0[8])) /* synthesis lut_function=(!(A)) */ ;
    defparam i4_1_lut.init = 16'h5555;
    LUT4 i6896_4_lut_4_lut (.A(n14083), .B(\mXs_0[24] ), .C(eX_0[3]), 
         .D(n70764), .Z(buf_x[390])) /* synthesis lut_function=(A (B+(C (D)))+!A !(B (C (D))+!B !(C (D)))) */ ;
    defparam i6896_4_lut_4_lut.init = 16'hbccc;
    LUT4 i18_3_lut_4_lut (.A(n14083), .B(\mXs_0[24] ), .C(eX_0[0]), .D(mXs_0[22]), 
         .Z(buf_x[111])) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam i18_3_lut_4_lut.init = 16'hfb0b;
    LUT4 buf_x_286__bdd_3_lut_4_lut (.A(n70807), .B(eX_0[2]), .C(n14083), 
         .D(\mXs_0[24] ), .Z(n69016)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (D)) */ ;
    defparam buf_x_286__bdd_3_lut_4_lut.init = 16'hf788;
    LUT4 i54637_else_3_lut (.A(buf_x[615]), .B(buf_r[38]), .C(eX_x[10]), 
         .Z(n70878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54637_else_3_lut.init = 16'hcaca;
    LUT4 i29132_2_lut (.A(eX_0[2]), .B(eX_0[3]), .Z(n40725)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i29132_2_lut.init = 16'heeee;
    LUT4 i67_4_lut (.A(mXs_0[0]), .B(buf_x[90]), .C(eX_0[1]), .D(eX_0[0]), 
         .Z(buf_x[178])) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;
    defparam i67_4_lut.init = 16'h0cac;
    LUT4 mux_14_i1_3_lut (.A(\exp_a[0] ), .B(n14059[0]), .C(\mXs_0[24] ), 
         .Z(mXs_0[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i1_3_lut.init = 16'hcaca;
    LUT4 i40_3_lut (.A(mXs_0[0]), .B(mXs_0[1]), .C(eX_0[0]), .Z(buf_x[89])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i40_3_lut.init = 16'hacac;
    LUT4 mux_14_i2_3_lut (.A(\exp_a[1] ), .B(n14059[1]), .C(\mXs_0[24] ), 
         .Z(mXs_0[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i2_3_lut.init = 16'hcaca;
    LUT4 i39_3_lut (.A(mXs_0[1]), .B(mXs_0[2]), .C(eX_0[0]), .Z(buf_x[90])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i39_3_lut.init = 16'hacac;
    LUT4 mux_14_i3_3_lut (.A(\exp_a[2] ), .B(n14059[2]), .C(\mXs_0[24] ), 
         .Z(mXs_0[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i3_3_lut.init = 16'hcaca;
    LUT4 i38_3_lut (.A(mXs_0[2]), .B(mXs_0[3]), .C(eX_0[0]), .Z(buf_x[91])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i38_3_lut.init = 16'hacac;
    LUT4 mux_14_i4_3_lut (.A(\exp_a[3] ), .B(n14059[3]), .C(\mXs_0[24] ), 
         .Z(mXs_0[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i4_3_lut.init = 16'hcaca;
    LUT4 i37_3_lut (.A(mXs_0[3]), .B(mXs_0[4]), .C(eX_0[0]), .Z(buf_x[92])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i37_3_lut.init = 16'hacac;
    LUT4 i54637_then_3_lut (.A(buf_r[6]), .B(buf_r[22]), .C(eX_x[10]), 
         .Z(n70879)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54637_then_3_lut.init = 16'hacac;
    LUT4 mux_14_i5_3_lut (.A(\exp_a[4] ), .B(n14059[4]), .C(\mXs_0[24] ), 
         .Z(mXs_0[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i5_3_lut.init = 16'hcaca;
    LUT4 i36_3_lut (.A(mXs_0[4]), .B(mXs_0[5]), .C(eX_0[0]), .Z(buf_x[93])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i36_3_lut.init = 16'hacac;
    LUT4 mux_14_i6_3_lut (.A(\exp_a[5] ), .B(n14059[5]), .C(\mXs_0[24] ), 
         .Z(mXs_0[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i6_3_lut.init = 16'hcaca;
    LUT4 i35_3_lut (.A(mXs_0[5]), .B(mXs_0[6]), .C(eX_0[0]), .Z(buf_x[94])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i35_3_lut.init = 16'hacac;
    LUT4 mux_14_i7_3_lut (.A(\exp_a[6] ), .B(n14059[6]), .C(\mXs_0[24] ), 
         .Z(mXs_0[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i7_3_lut.init = 16'hcaca;
    LUT4 i34_3_lut (.A(mXs_0[6]), .B(mXs_0[7]), .C(eX_0[0]), .Z(buf_x[95])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i34_3_lut.init = 16'hacac;
    LUT4 mux_14_i8_3_lut (.A(\exp_a[7] ), .B(n14059[7]), .C(\mXs_0[24] ), 
         .Z(mXs_0[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i8_3_lut.init = 16'hcaca;
    LUT4 i33_3_lut (.A(mXs_0[7]), .B(mXs_0[8]), .C(eX_0[0]), .Z(buf_x[96])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i33_3_lut.init = 16'hacac;
    LUT4 mux_14_i9_3_lut (.A(\exp_a[8] ), .B(n14059[8]), .C(\mXs_0[24] ), 
         .Z(mXs_0[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i9_3_lut.init = 16'hcaca;
    LUT4 i32_3_lut (.A(mXs_0[8]), .B(mXs_0[9]), .C(eX_0[0]), .Z(buf_x[97])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i32_3_lut.init = 16'hacac;
    LUT4 mux_14_i10_3_lut (.A(\exp_a[9] ), .B(n14059[9]), .C(\mXs_0[24] ), 
         .Z(mXs_0[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i10_3_lut.init = 16'hcaca;
    LUT4 i31_3_lut (.A(mXs_0[9]), .B(mXs_0[10]), .C(eX_0[0]), .Z(buf_x[98])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i31_3_lut.init = 16'hacac;
    LUT4 mux_14_i11_3_lut (.A(\exp_a[10] ), .B(n14059[10]), .C(\mXs_0[24] ), 
         .Z(mXs_0[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i11_3_lut.init = 16'hcaca;
    LUT4 i30_3_lut (.A(mXs_0[10]), .B(mXs_0[11]), .C(eX_0[0]), .Z(buf_x[99])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i30_3_lut.init = 16'hacac;
    LUT4 mux_14_i12_3_lut (.A(\exp_a[11] ), .B(n14059[11]), .C(\mXs_0[24] ), 
         .Z(mXs_0[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i12_3_lut.init = 16'hcaca;
    LUT4 i29_3_lut (.A(mXs_0[11]), .B(mXs_0[12]), .C(eX_0[0]), .Z(buf_x[100])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i29_3_lut.init = 16'hacac;
    LUT4 mux_14_i13_3_lut (.A(\exp_a[12] ), .B(n14059[12]), .C(\mXs_0[24] ), 
         .Z(mXs_0[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i13_3_lut.init = 16'hcaca;
    LUT4 i28_3_lut (.A(mXs_0[12]), .B(mXs_0[13]), .C(eX_0[0]), .Z(buf_x[101])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i28_3_lut.init = 16'hacac;
    LUT4 mux_14_i14_3_lut (.A(\exp_a[13] ), .B(n14059[13]), .C(\mXs_0[24] ), 
         .Z(mXs_0[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i14_3_lut.init = 16'hcaca;
    LUT4 i27_3_lut (.A(mXs_0[13]), .B(mXs_0[14]), .C(eX_0[0]), .Z(buf_x[102])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i27_3_lut.init = 16'hacac;
    LUT4 mux_14_i15_3_lut (.A(\exp_a[14] ), .B(n14059[14]), .C(\mXs_0[24] ), 
         .Z(mXs_0[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i15_3_lut.init = 16'hcaca;
    LUT4 i26_3_lut (.A(mXs_0[14]), .B(mXs_0[15]), .C(eX_0[0]), .Z(buf_x[103])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i26_3_lut.init = 16'hacac;
    LUT4 mux_14_i16_3_lut (.A(\exp_a[15] ), .B(n14059[15]), .C(\mXs_0[24] ), 
         .Z(mXs_0[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i16_3_lut.init = 16'hcaca;
    LUT4 i25_3_lut (.A(mXs_0[15]), .B(mXs_0[16]), .C(eX_0[0]), .Z(buf_x[104])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i25_3_lut.init = 16'hacac;
    LUT4 mux_14_i17_3_lut (.A(\exp_a[16] ), .B(n14059[16]), .C(\mXs_0[24] ), 
         .Z(mXs_0[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i17_3_lut.init = 16'hcaca;
    LUT4 i24_3_lut (.A(mXs_0[16]), .B(mXs_0[17]), .C(eX_0[0]), .Z(buf_x[105])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i24_3_lut.init = 16'hacac;
    LUT4 i110_3_lut (.A(buf_x[287]), .B(\mXs_0[24] ), .C(eX_0[3]), .Z(buf_x[383])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i110_3_lut.init = 16'hacac;
    LUT4 mux_14_i18_3_lut (.A(\exp_a[17] ), .B(n14059[17]), .C(\mXs_0[24] ), 
         .Z(mXs_0[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i18_3_lut.init = 16'hcaca;
    LUT4 i23_3_lut (.A(mXs_0[17]), .B(mXs_0[18]), .C(eX_0[0]), .Z(buf_x[106])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i23_3_lut.init = 16'hacac;
    LUT4 i109_3_lut (.A(buf_x[288]), .B(\mXs_0[24] ), .C(eX_0[3]), .Z(buf_x[384])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i109_3_lut.init = 16'hacac;
    LUT4 mux_14_i19_3_lut (.A(\exp_a[18] ), .B(n14059[18]), .C(\mXs_0[24] ), 
         .Z(mXs_0[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i19_3_lut.init = 16'hcaca;
    LUT4 i22_3_lut (.A(mXs_0[18]), .B(mXs_0[19]), .C(eX_0[0]), .Z(buf_x[107])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i22_3_lut.init = 16'hacac;
    LUT4 i108_3_lut (.A(buf_x[289]), .B(\mXs_0[24] ), .C(eX_0[3]), .Z(buf_x[385])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i108_3_lut.init = 16'hacac;
    LUT4 mux_14_i20_3_lut (.A(\exp_a[19] ), .B(n14059[19]), .C(\mXs_0[24] ), 
         .Z(mXs_0[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i20_3_lut.init = 16'hcaca;
    LUT4 i21_3_lut (.A(mXs_0[19]), .B(mXs_0[20]), .C(eX_0[0]), .Z(buf_x[108])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i21_3_lut.init = 16'hacac;
    LUT4 i107_3_lut (.A(buf_x[290]), .B(\mXs_0[24] ), .C(eX_0[3]), .Z(buf_x[386])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i107_3_lut.init = 16'hacac;
    LUT4 mux_14_i21_3_lut (.A(\exp_a[20] ), .B(n14059[20]), .C(\mXs_0[24] ), 
         .Z(mXs_0[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i21_3_lut.init = 16'hcaca;
    LUT4 i20_3_lut (.A(mXs_0[20]), .B(mXs_0[21]), .C(eX_0[0]), .Z(buf_x[109])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i20_3_lut.init = 16'hacac;
    LUT4 mux_14_i22_3_lut (.A(\exp_a[21] ), .B(n14059[21]), .C(\mXs_0[24] ), 
         .Z(mXs_0[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i22_3_lut.init = 16'hcaca;
    LUT4 i19_3_lut (.A(mXs_0[21]), .B(mXs_0[22]), .C(eX_0[0]), .Z(buf_x[110])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i19_3_lut.init = 16'hacac;
    LUT4 mux_14_i23_3_lut (.A(\exp_a[22] ), .B(n14059[22]), .C(\mXs_0[24] ), 
         .Z(mXs_0[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_14_i23_3_lut.init = 16'hcaca;
    LUT4 i6898_4_lut (.A(\mXs_0[24] ), .B(buf_x[111]), .C(n70806), .D(eX_0[3]), 
         .Z(buf_x[389])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6898_4_lut.init = 16'hcaaa;
    PFUMX i56080 (.BLUT(n70875), .ALUT(n70876), .C0(\eX_x[11] ), .Z(\nX_a0[30] ));
    LUT4 i216_3_lut (.A(buf_r[7]), .B(buf_r[23]), .C(eX_x[10]), .Z(\buf_x[463] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i216_3_lut.init = 16'hacac;
    FD1S3IX buf_r_0__367 (.D(mXs_0[0]), .CK(clock), .CD(n41668), .Q(buf_r[0]));
    defparam buf_r_0__367.GSR = "DISABLED";
    FD1S3IX buf_r_1__366 (.D(buf_x[89]), .CK(clock), .CD(n41530), .Q(buf_r[1]));
    defparam buf_r_1__366.GSR = "DISABLED";
    FD1S3IX buf_r_3__364 (.D(buf_x[179]), .CK(clock), .CD(n40725), .Q(buf_r[3]));
    defparam buf_r_3__364.GSR = "DISABLED";
    LUT4 i54634_else_3_lut (.A(buf_x[615]), .B(buf_r[37]), .C(eX_x[10]), 
         .Z(n70875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54634_else_3_lut.init = 16'hcaca;
    LUT4 buf_x_110__bdd_3_lut (.A(eX_0[0]), .B(\mXs_0[24] ), .C(n14083), 
         .Z(n69147)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;
    defparam buf_x_110__bdd_3_lut.init = 16'he6e6;
    PFUMX i55441 (.BLUT(n69147), .ALUT(buf_x[110]), .C0(eX_0[1]), .Z(buf_x[200]));
    LUT4 i54634_then_3_lut (.A(buf_r[5]), .B(buf_r[21]), .C(eX_x[10]), 
         .Z(n70876)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54634_then_3_lut.init = 16'hacac;
    CCU2D add_4_9 (.A0(\exp_a[30] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61695), 
          .S1(n4));
    defparam add_4_9.INIT0 = 16'h5555;
    defparam add_4_9.INIT1 = 16'h0000;
    defparam add_4_9.INJECT1_0 = "NO";
    defparam add_4_9.INJECT1_1 = "NO";
    CCU2D add_4_7 (.A0(\exp_a[28] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[29] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61694), .COUT(n61695), .S0(eX_0[5]));
    defparam add_4_7.INIT0 = 16'h5aaa;
    defparam add_4_7.INIT1 = 16'h5aaa;
    defparam add_4_7.INJECT1_0 = "NO";
    defparam add_4_7.INJECT1_1 = "NO";
    CCU2D add_4_5 (.A0(\exp_a[26] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[27] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61693), .COUT(n61694), .S0(eX_0[3]), .S1(eX_0[4]));
    defparam add_4_5.INIT0 = 16'h5555;
    defparam add_4_5.INIT1 = 16'h5555;
    defparam add_4_5.INJECT1_0 = "NO";
    defparam add_4_5.INJECT1_1 = "NO";
    PFUMX i55408 (.BLUT(n69079), .ALUT(buf_x[198]), .C0(eX_0[2]), .Z(buf_x[290]));
    CCU2D add_4_3 (.A0(\exp_a[24] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[25] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61692), .COUT(n61693), .S0(eX_0[1]), .S1(eX_0[2]));
    defparam add_4_3.INIT0 = 16'h5aaa;
    defparam add_4_3.INIT1 = 16'h5555;
    defparam add_4_3.INJECT1_0 = "NO";
    defparam add_4_3.INJECT1_1 = "NO";
    CCU2D add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[23] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n61692), .S1(eX_0[0]));
    defparam add_4_1.INIT0 = 16'hF000;
    defparam add_4_1.INIT1 = 16'h5555;
    defparam add_4_1.INJECT1_0 = "NO";
    defparam add_4_1.INJECT1_1 = "NO";
    LUT4 i212_3_lut (.A(buf_r[11]), .B(buf_r[27]), .C(eX_x[10]), .Z(\buf_x[467] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i212_3_lut.init = 16'hacac;
    LUT4 i211_3_lut (.A(buf_r[12]), .B(buf_r[28]), .C(eX_x[10]), .Z(\buf_x[468] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i211_3_lut.init = 16'hacac;
    LUT4 i210_3_lut (.A(buf_r[13]), .B(buf_r[29]), .C(eX_x[10]), .Z(\buf_x[469] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i210_3_lut.init = 16'hacac;
    LUT4 i209_3_lut (.A(buf_r[14]), .B(buf_r[30]), .C(eX_x[10]), .Z(\buf_x[470] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i209_3_lut.init = 16'hacac;
    LUT4 i208_3_lut (.A(buf_r[15]), .B(buf_r[31]), .C(eX_x[10]), .Z(\buf_x[471] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i208_3_lut.init = 16'hacac;
    LUT4 i272_3_lut (.A(\buf_x[463] ), .B(buf_x[615]), .C(\eX_x[11] ), 
         .Z(\nX_a0[32] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i272_3_lut.init = 16'hacac;
    LUT4 i215_3_lut (.A(buf_r[8]), .B(buf_r[24]), .C(eX_x[10]), .Z(\buf_x[464] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i215_3_lut.init = 16'hacac;
    LUT4 i271_3_lut (.A(\buf_x[464] ), .B(buf_x[615]), .C(\eX_x[11] ), 
         .Z(\nX_a0[33] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i271_3_lut.init = 16'hacac;
    LUT4 i214_3_lut (.A(buf_r[9]), .B(buf_r[25]), .C(eX_x[10]), .Z(\buf_x[465] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i214_3_lut.init = 16'hacac;
    LUT4 i270_3_lut (.A(\buf_x[465] ), .B(buf_x[615]), .C(\eX_x[11] ), 
         .Z(\nX_a0[34] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i270_3_lut.init = 16'hacac;
    LUT4 i213_3_lut (.A(buf_r[10]), .B(buf_r[26]), .C(eX_x[10]), .Z(\buf_x[466] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i213_3_lut.init = 16'hacac;
    LUT4 i269_3_lut (.A(\buf_x[466] ), .B(buf_x[615]), .C(\eX_x[11] ), 
         .Z(\nX_a0[35] )) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i269_3_lut.init = 16'hacac;
    PFUMX i55375 (.BLUT(n69021), .ALUT(buf_x[197]), .C0(eX_0[2]), .Z(buf_x[289]));
    LUT4 buf_x_197__bdd_3_lut (.A(buf_x[111]), .B(eX_0[1]), .C(\mXs_0[24] ), 
         .Z(n69021)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam buf_x_197__bdd_3_lut.init = 16'hb8b8;
    PFUMX i55371 (.BLUT(n69016), .ALUT(buf_x[286]), .C0(eX_0[3]), .Z(buf_x[382]));
    PFUMX i55369 (.BLUT(n69010), .ALUT(buf_x[285]), .C0(eX_0[3]), .Z(buf_x[381]));
    PFUMX i55367 (.BLUT(n69008), .ALUT(buf_x[284]), .C0(eX_0[3]), .Z(buf_x[380]));
    LUT4 buf_x_284__bdd_3_lut (.A(buf_x[200]), .B(eX_0[2]), .C(\mXs_0[24] ), 
         .Z(n69008)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam buf_x_284__bdd_3_lut.init = 16'hb8b8;
    PFUMX i55365 (.BLUT(n69004), .ALUT(buf_x[283]), .C0(eX_0[3]), .Z(buf_x[379]));
    LUT4 buf_x_283__bdd_3_lut (.A(buf_x[199]), .B(eX_0[2]), .C(\mXs_0[24] ), 
         .Z(n69004)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam buf_x_283__bdd_3_lut.init = 16'hb8b8;
    PFUMX i56126 (.BLUT(n70944), .ALUT(n70945), .C0(eX_x[10]), .Z(\nX_a0[24] ));
    LUT4 i280_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[15]), 
         .Z(n70944)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i280_else_2_lut.init = 16'he2e2;
    LUT4 i280_then_2_lut (.A(buf_r[31]), .B(\eX_x[11] ), .Z(n70945)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i280_then_2_lut.init = 16'h2222;
    PFUMX i56124 (.BLUT(n70941), .ALUT(n70942), .C0(eX_x[10]), .Z(\nX_a0[23] ));
    LUT4 i281_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[14]), 
         .Z(n70941)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i281_else_2_lut.init = 16'he2e2;
    LUT4 i281_then_2_lut (.A(buf_r[30]), .B(\eX_x[11] ), .Z(n70942)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i281_then_2_lut.init = 16'h2222;
    PFUMX i56122 (.BLUT(n70938), .ALUT(n70939), .C0(eX_x[10]), .Z(\nX_a0[22] ));
    LUT4 i282_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[13]), 
         .Z(n70938)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i282_else_2_lut.init = 16'he2e2;
    LUT4 i282_then_2_lut (.A(buf_r[29]), .B(\eX_x[11] ), .Z(n70939)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i282_then_2_lut.init = 16'h2222;
    PFUMX i56120 (.BLUT(n70935), .ALUT(n70936), .C0(eX_x[10]), .Z(\nX_a0[21] ));
    LUT4 i283_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[12]), 
         .Z(n70935)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i283_else_2_lut.init = 16'he2e2;
    LUT4 i283_then_2_lut (.A(buf_r[28]), .B(\eX_x[11] ), .Z(n70936)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i283_then_2_lut.init = 16'h2222;
    CCU2D add_4598_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61634), 
          .S0(n14083));
    defparam add_4598_cout.INIT0 = 16'h0000;
    defparam add_4598_cout.INIT1 = 16'h0000;
    defparam add_4598_cout.INJECT1_0 = "NO";
    defparam add_4598_cout.INJECT1_1 = "NO";
    PFUMX i56118 (.BLUT(n70932), .ALUT(n70933), .C0(eX_x[10]), .Z(\nX_a0[20] ));
    LUT4 i284_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[11]), 
         .Z(n70932)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i284_else_2_lut.init = 16'he2e2;
    LUT4 i284_then_2_lut (.A(buf_r[27]), .B(\eX_x[11] ), .Z(n70933)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i284_then_2_lut.init = 16'h2222;
    CCU2D add_4598_23 (.A0(\exp_a[21] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[22] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61633), .COUT(n61634), .S0(n14059[21]), .S1(n14059[22]));
    defparam add_4598_23.INIT0 = 16'hf555;
    defparam add_4598_23.INIT1 = 16'hf555;
    defparam add_4598_23.INJECT1_0 = "NO";
    defparam add_4598_23.INJECT1_1 = "NO";
    CCU2D add_4598_21 (.A0(\exp_a[19] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[20] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61632), .COUT(n61633), .S0(n14059[19]), .S1(n14059[20]));
    defparam add_4598_21.INIT0 = 16'hf555;
    defparam add_4598_21.INIT1 = 16'hf555;
    defparam add_4598_21.INJECT1_0 = "NO";
    defparam add_4598_21.INJECT1_1 = "NO";
    PFUMX i56116 (.BLUT(n70929), .ALUT(n70930), .C0(eX_x[10]), .Z(\nX_a0[19] ));
    LUT4 i285_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[10]), 
         .Z(n70929)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i285_else_2_lut.init = 16'he2e2;
    LUT4 i285_then_2_lut (.A(buf_r[26]), .B(\eX_x[11] ), .Z(n70930)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i285_then_2_lut.init = 16'h2222;
    PFUMX i56114 (.BLUT(n70926), .ALUT(n70927), .C0(eX_x[10]), .Z(\nX_a0[18] ));
    LUT4 i286_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[9]), 
         .Z(n70926)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i286_else_2_lut.init = 16'he2e2;
    LUT4 i286_then_2_lut (.A(buf_r[25]), .B(\eX_x[11] ), .Z(n70927)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i286_then_2_lut.init = 16'h2222;
    CCU2D add_4598_19 (.A0(\exp_a[17] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[18] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61631), .COUT(n61632), .S0(n14059[17]), .S1(n14059[18]));
    defparam add_4598_19.INIT0 = 16'hf555;
    defparam add_4598_19.INIT1 = 16'hf555;
    defparam add_4598_19.INJECT1_0 = "NO";
    defparam add_4598_19.INJECT1_1 = "NO";
    CCU2D add_4598_17 (.A0(\exp_a[15] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[16] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61630), .COUT(n61631), .S0(n14059[15]), .S1(n14059[16]));
    defparam add_4598_17.INIT0 = 16'hf555;
    defparam add_4598_17.INIT1 = 16'hf555;
    defparam add_4598_17.INJECT1_0 = "NO";
    defparam add_4598_17.INJECT1_1 = "NO";
    CCU2D add_4598_15 (.A0(\exp_a[13] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61629), .COUT(n61630), .S0(n14059[13]), .S1(n14059[14]));
    defparam add_4598_15.INIT0 = 16'hf555;
    defparam add_4598_15.INIT1 = 16'hf555;
    defparam add_4598_15.INJECT1_0 = "NO";
    defparam add_4598_15.INJECT1_1 = "NO";
    PFUMX i56110 (.BLUT(n70920), .ALUT(n70921), .C0(eX_x[10]), .Z(\nX_a0[17] ));
    LUT4 i287_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[8]), 
         .Z(n70920)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i287_else_2_lut.init = 16'he2e2;
    LUT4 i287_then_2_lut (.A(buf_r[24]), .B(\eX_x[11] ), .Z(n70921)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i287_then_2_lut.init = 16'h2222;
    CCU2D add_4598_13 (.A0(\exp_a[11] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[12] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61628), .COUT(n61629), .S0(n14059[11]), .S1(n14059[12]));
    defparam add_4598_13.INIT0 = 16'hf555;
    defparam add_4598_13.INIT1 = 16'hf555;
    defparam add_4598_13.INJECT1_0 = "NO";
    defparam add_4598_13.INJECT1_1 = "NO";
    PFUMX i56108 (.BLUT(n70917), .ALUT(n70918), .C0(eX_x[10]), .Z(\nX_a0[16] ));
    CCU2D add_4598_11 (.A0(\exp_a[9] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[10] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61627), .COUT(n61628), .S0(n14059[9]), .S1(n14059[10]));
    defparam add_4598_11.INIT0 = 16'hf555;
    defparam add_4598_11.INIT1 = 16'hf555;
    defparam add_4598_11.INJECT1_0 = "NO";
    defparam add_4598_11.INJECT1_1 = "NO";
    CCU2D add_4598_9 (.A0(\exp_a[7] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[8] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61626), .COUT(n61627), .S0(n14059[7]), .S1(n14059[8]));
    defparam add_4598_9.INIT0 = 16'hf555;
    defparam add_4598_9.INIT1 = 16'hf555;
    defparam add_4598_9.INJECT1_0 = "NO";
    defparam add_4598_9.INJECT1_1 = "NO";
    LUT4 i288_else_2_lut (.A(buf_x[615]), .B(\eX_x[11] ), .C(buf_r[7]), 
         .Z(n70917)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i288_else_2_lut.init = 16'he2e2;
    LUT4 i288_then_2_lut (.A(buf_r[23]), .B(\eX_x[11] ), .Z(n70918)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i288_then_2_lut.init = 16'h2222;
    PFUMX i56106 (.BLUT(n70914), .ALUT(n70915), .C0(\eX_x[11] ), .Z(\nX_a0[15] ));
    LUT4 i23137_else_2_lut (.A(buf_r[38]), .B(eX_x[10]), .C(buf_r[22]), 
         .Z(n70914)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23137_else_2_lut.init = 16'he2e2;
    LUT4 i23137_then_2_lut (.A(buf_r[6]), .B(eX_x[10]), .Z(n70915)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23137_then_2_lut.init = 16'h2222;
    PFUMX i56104 (.BLUT(n70911), .ALUT(n70912), .C0(\eX_x[11] ), .Z(\nX_a0[14] ));
    LUT4 i23148_else_2_lut (.A(buf_r[37]), .B(eX_x[10]), .C(buf_r[21]), 
         .Z(n70911)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23148_else_2_lut.init = 16'he2e2;
    LUT4 i23148_then_2_lut (.A(buf_r[5]), .B(eX_x[10]), .Z(n70912)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23148_then_2_lut.init = 16'h2222;
    PFUMX i56102 (.BLUT(n70908), .ALUT(n70909), .C0(\eX_x[11] ), .Z(\nX_a0[13] ));
    LUT4 i23159_else_2_lut (.A(buf_r[36]), .B(eX_x[10]), .C(buf_r[20]), 
         .Z(n70908)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23159_else_2_lut.init = 16'he2e2;
    LUT4 i23159_then_2_lut (.A(buf_r[4]), .B(eX_x[10]), .Z(n70909)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23159_then_2_lut.init = 16'h2222;
    PFUMX i56100 (.BLUT(n70905), .ALUT(n70906), .C0(\eX_x[11] ), .Z(\nX_a0[12] ));
    LUT4 i23170_else_2_lut (.A(buf_r[35]), .B(eX_x[10]), .C(buf_r[19]), 
         .Z(n70905)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23170_else_2_lut.init = 16'he2e2;
    LUT4 i23170_then_2_lut (.A(buf_r[3]), .B(eX_x[10]), .Z(n70906)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23170_then_2_lut.init = 16'h2222;
    PFUMX i56098 (.BLUT(n70902), .ALUT(n70903), .C0(\eX_x[11] ), .Z(\nX_a0[11] ));
    CCU2D add_4598_7 (.A0(\exp_a[5] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[6] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61625), .COUT(n61626), .S0(n14059[5]), .S1(n14059[6]));
    defparam add_4598_7.INIT0 = 16'hf555;
    defparam add_4598_7.INIT1 = 16'hf555;
    defparam add_4598_7.INJECT1_0 = "NO";
    defparam add_4598_7.INJECT1_1 = "NO";
    LUT4 i23181_else_2_lut (.A(buf_r[34]), .B(eX_x[10]), .C(buf_r[18]), 
         .Z(n70902)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23181_else_2_lut.init = 16'he2e2;
    LUT4 i23181_then_2_lut (.A(buf_r[2]), .B(eX_x[10]), .Z(n70903)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23181_then_2_lut.init = 16'h2222;
    CCU2D add_4598_5 (.A0(\exp_a[3] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[4] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61624), .COUT(n61625), .S0(n14059[3]), .S1(n14059[4]));
    defparam add_4598_5.INIT0 = 16'hf555;
    defparam add_4598_5.INIT1 = 16'hf555;
    defparam add_4598_5.INJECT1_0 = "NO";
    defparam add_4598_5.INJECT1_1 = "NO";
    CCU2D add_4598_3 (.A0(\exp_a[1] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[2] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61623), .COUT(n61624), .S0(n14059[1]), .S1(n14059[2]));
    defparam add_4598_3.INIT0 = 16'hf555;
    defparam add_4598_3.INIT1 = 16'hf555;
    defparam add_4598_3.INJECT1_0 = "NO";
    defparam add_4598_3.INJECT1_1 = "NO";
    CCU2D add_4598_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\exp_a[0] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n61623), .S1(n14059[0]));
    defparam add_4598_1.INIT0 = 16'hF000;
    defparam add_4598_1.INIT1 = 16'h0aaa;
    defparam add_4598_1.INJECT1_0 = "NO";
    defparam add_4598_1.INJECT1_1 = "NO";
    PFUMX i56096 (.BLUT(n70899), .ALUT(n70900), .C0(\eX_x[11] ), .Z(\nX_a0[10] ));
    LUT4 i23192_else_2_lut (.A(buf_r[33]), .B(eX_x[10]), .C(buf_r[17]), 
         .Z(n70899)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23192_else_2_lut.init = 16'he2e2;
    LUT4 i23192_then_2_lut (.A(buf_r[1]), .B(eX_x[10]), .Z(n70900)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23192_then_2_lut.init = 16'h2222;
    PFUMX i56094 (.BLUT(n70896), .ALUT(n70897), .C0(\eX_x[11] ), .Z(\nX_a0[9] ));
    LUT4 i23203_else_2_lut (.A(buf_r[32]), .B(eX_x[10]), .C(buf_r[16]), 
         .Z(n70896)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam i23203_else_2_lut.init = 16'he2e2;
    LUT4 i23203_then_2_lut (.A(buf_r[0]), .B(eX_x[10]), .Z(n70897)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i23203_then_2_lut.init = 16'h2222;
    PFUMX i56092 (.BLUT(n70893), .ALUT(n70894), .C0(\eX_x[11] ), .Z(\nX_a0[25] ));
    LUT4 i54652_else_3_lut (.A(buf_x[615]), .B(buf_r[32]), .C(eX_x[10]), 
         .Z(n70893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54652_else_3_lut.init = 16'hcaca;
    LUT4 i54652_then_3_lut (.A(buf_r[0]), .B(buf_r[16]), .C(eX_x[10]), 
         .Z(n70894)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54652_then_3_lut.init = 16'hacac;
    PFUMX i56090 (.BLUT(n70890), .ALUT(n70891), .C0(\eX_x[11] ), .Z(\nX_a0[26] ));
    LUT4 i54649_else_3_lut (.A(buf_x[615]), .B(buf_r[33]), .C(eX_x[10]), 
         .Z(n70890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54649_else_3_lut.init = 16'hcaca;
    LUT4 i54649_then_3_lut (.A(buf_r[1]), .B(buf_r[17]), .C(eX_x[10]), 
         .Z(n70891)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54649_then_3_lut.init = 16'hacac;
    PFUMX i56088 (.BLUT(n70887), .ALUT(n70888), .C0(\eX_x[11] ), .Z(\nX_a0[27] ));
    LUT4 i54646_else_3_lut (.A(buf_x[615]), .B(buf_r[34]), .C(eX_x[10]), 
         .Z(n70887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54646_else_3_lut.init = 16'hcaca;
    LUT4 i54646_then_3_lut (.A(buf_r[2]), .B(buf_r[18]), .C(eX_x[10]), 
         .Z(n70888)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54646_then_3_lut.init = 16'hacac;
    PFUMX i56086 (.BLUT(n70884), .ALUT(n70885), .C0(\eX_x[11] ), .Z(\nX_a0[28] ));
    LUT4 i54643_else_3_lut (.A(buf_x[615]), .B(buf_r[35]), .C(eX_x[10]), 
         .Z(n70884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54643_else_3_lut.init = 16'hcaca;
    LUT4 i54643_then_3_lut (.A(buf_r[3]), .B(buf_r[19]), .C(eX_x[10]), 
         .Z(n70885)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i54643_then_3_lut.init = 16'hacac;
    PFUMX i56084 (.BLUT(n70881), .ALUT(n70882), .C0(\eX_x[11] ), .Z(\nX_a0[29] ));
    \delay(1,1)  delay_ufl (.nX_d({nX_d}), .clock(clock), .\eX_0[8] (eX_0[8]));
    
endmodule
//
// Verilog Description of module \delay(1,1) 
//

module \delay(1,1)  (nX_d, clock, \eX_0[8] );
    output [0:0]nX_d;
    input clock;
    input \eX_0[8] ;
    
    
    FD1S3AX buf_1__5 (.D(\eX_0[8] ), .CK(clock), .Q(nX_d[0]));
    defparam buf_1__5.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \mult_clk(28,22,false,false,0,2) 
//

module \mult_clk(28,22,false,false,0,2)  (nEY1_d2, nZ0_d2, GND_net, clock, 
            n23965, n23964, n23963, n23962, n23961, n23960, n23959, 
            n23958, n23957, n23956, \nZ1_e0[48] , \nZ1_e0[49] , \nZ1_e0[46] , 
            \nZ1_e0[47] , \nZ1_e0[44] , \nZ1_e0[45] , \nZ1_e0[42] , 
            \nZ1_e0[43] , \nZ1_e0[40] , \nZ1_e0[41] , \nZ1_e0[38] , 
            \nZ1_e0[39] , \nZ1_e0[36] , \nZ1_e0[37] , \nZ1_e0[34] , 
            \nZ1_e0[35] , \nZ1_e0[32] , \nZ1_e0[33] , \nZ1_e0[30] , 
            \nZ1_e0[31] , \nZ1_e0[29] );
    input [27:0]nEY1_d2;
    input [21:0]nZ0_d2;
    input GND_net;
    input clock;
    input n23965;
    input n23964;
    input n23963;
    input n23962;
    input n23961;
    input n23960;
    input n23959;
    input n23958;
    input n23957;
    input n23956;
    output \nZ1_e0[48] ;
    output \nZ1_e0[49] ;
    output \nZ1_e0[46] ;
    output \nZ1_e0[47] ;
    output \nZ1_e0[44] ;
    output \nZ1_e0[45] ;
    output \nZ1_e0[42] ;
    output \nZ1_e0[43] ;
    output \nZ1_e0[40] ;
    output \nZ1_e0[41] ;
    output \nZ1_e0[38] ;
    output \nZ1_e0[39] ;
    output \nZ1_e0[36] ;
    output \nZ1_e0[37] ;
    output \nZ1_e0[34] ;
    output \nZ1_e0[35] ;
    output \nZ1_e0[32] ;
    output \nZ1_e0[33] ;
    output \nZ1_e0[30] ;
    output \nZ1_e0[31] ;
    output \nZ1_e0[29] ;
    
    wire [2018:0]buf_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [2018:0]buf_r;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(337[10:15])
    
    wire n61975, n61976, n61974, n61973, n61972, n61971, n61970, 
        n61969, n61968, n61967, n61966, n61965, n61964, n61963, 
        n61962, n61961, n61960, n61959, n61958, n61957, n61956, 
        n61955, n61954, n61953, n61952, n61951, n61950, n61949, 
        n61948, n61947, n61946, n61945, n61944, n61943, n61942, 
        n61941, n61940, n61939, n61938, n61937, n61936, n61935, 
        n61934, n61933, n61932, n61931, n61930, n61929, n61928, 
        n61927, n61926, n61925, n61924, n61923, n61922, n61921, 
        n61920, n61919, n61918, n61917, n61916, n61915, n61914, 
        n61913, n61912, n61911, n61910, n61909, n61908, n61907, 
        n61906, n61905, n61904, n61903, n61902, n61901, n61900, 
        n61899, n61898, n61897, n61896, n61895, n61894, n61893, 
        n61892, n61891, n61890, n61889, n61888, n61887, n61886, 
        n61885, n61884, n61883, n61882, n61881, n61880, n61879, 
        n61878, n61877, n61876, n61875, n61874, n61873, n61872, 
        n61871, n61870, n61869, n61868, n61867, n61866, n61865, 
        n61864, n61863, n61862, n61861, n61854, n61853, n61852, 
        n61851, n61850, n61849, n61848, n61847, n61846, n61845, 
        n61844, n61843, n61842, n61841, n61779, n61778, n61777, 
        n61776, n61775, n61774, n61773, n61772, n61771, n61770, 
        n61769, n61768, n61767, n61766, n62154, n62153, n62152, 
        n62151, n62150, n62149, n62148, n62147, n62146, n62145, 
        n62144, n62143, n62142, n62141, n62140, n62139, n62138, 
        n62137, n62136, n62135, n62134, n62133, n62132, n62131, 
        n62130, n62129, n62128, n62127, n62126, n62125, n62124, 
        n62123, n62122, n62121, n62116, n62115, n62114, n62113, 
        n62112, n62111, n62110, n62109, n62108, n62107, n62106, 
        n62105, n62104, n62103, n62102, n62101, n62099, n62098, 
        n62097, n62096, n62095, n62094, n62093, n62092, n62091, 
        n62090, n62089, n62088, n62087, n62086, n62085, n62084, 
        n62079, n62078, n62077, n62076, n62075, n62074, n62073, 
        n62072, n62071, n62070, n62069, n62068, n62067, n62066, 
        n62065, n62063, n62062, n62061, n62060, n62059, n62058, 
        n62057, n62056, n62055, n62054, n62053, n62052, n62051, 
        n62050, n62049, n62047, n62046, n62045, n62044, n62043, 
        n62042, n62041, n62040, n62039, n62038, n62037, n62036, 
        n62035, n62034, n62033, n62031, n62030, n62029, n62028, 
        n62027, n62026, n62025, n62024, n62023, n62022, n62021, 
        n62020, n62019, n62018, n62017, n62015, n62014, n62013, 
        n62012, n62011, n62010, n62009, n62008, n62007, n62006, 
        n62005, n62004, n62003, n62002, n62001, n62000, n61999, 
        n61998, n61997, n61996, n61995, n61994, n61993, n61992, 
        n61991, n61990, n61989, n61988, n61987, n61986, n61985, 
        n61984, n61983, n61982, n61981, n61980, n61979, n61978, 
        n61977;
    
    CCU2D add_4612_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[18]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[7]), .B1(nZ0_d2[18]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[19]), .CIN(n61975), .COUT(n61976), .S0(buf_x[1245]), 
          .S1(buf_x[1246]));
    defparam add_4612_7.INIT0 = 16'h7888;
    defparam add_4612_7.INIT1 = 16'h7888;
    defparam add_4612_7.INJECT1_0 = "NO";
    defparam add_4612_7.INJECT1_1 = "NO";
    CCU2D add_4612_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[18]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[5]), .B1(nZ0_d2[18]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[19]), .CIN(n61974), .COUT(n61975), .S0(buf_x[1243]), 
          .S1(buf_x[1244]));
    defparam add_4612_5.INIT0 = 16'h7888;
    defparam add_4612_5.INIT1 = 16'h7888;
    defparam add_4612_5.INJECT1_0 = "NO";
    defparam add_4612_5.INJECT1_1 = "NO";
    CCU2D add_4612_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[18]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[3]), .B1(nZ0_d2[18]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[19]), .CIN(n61973), .COUT(n61974), .S0(buf_x[1241]), 
          .S1(buf_x[1242]));
    defparam add_4612_3.INIT0 = 16'h7888;
    defparam add_4612_3.INIT1 = 16'h7888;
    defparam add_4612_3.INJECT1_0 = "NO";
    defparam add_4612_3.INJECT1_1 = "NO";
    CCU2D add_4612_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[18]), .C1(nEY1_d2[0]), .D1(nZ0_d2[19]), 
          .COUT(n61973), .S1(buf_x[1240]));
    defparam add_4612_1.INIT0 = 16'hF000;
    defparam add_4612_1.INIT1 = 16'h7888;
    defparam add_4612_1.INJECT1_0 = "NO";
    defparam add_4612_1.INJECT1_1 = "NO";
    CCU2D add_4611_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[17]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61972), .S0(buf_x[1236]), .S1(buf_x[1237]));
    defparam add_4611_29.INIT0 = 16'h7888;
    defparam add_4611_29.INIT1 = 16'h0000;
    defparam add_4611_29.INJECT1_0 = "NO";
    defparam add_4611_29.INJECT1_1 = "NO";
    CCU2D add_4611_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[16]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[27]), .B1(nZ0_d2[16]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[17]), .CIN(n61971), .COUT(n61972), .S0(buf_x[1234]), 
          .S1(buf_x[1235]));
    defparam add_4611_27.INIT0 = 16'h7888;
    defparam add_4611_27.INIT1 = 16'h7888;
    defparam add_4611_27.INJECT1_0 = "NO";
    defparam add_4611_27.INJECT1_1 = "NO";
    CCU2D add_4611_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[16]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[25]), .B1(nZ0_d2[16]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[17]), .CIN(n61970), .COUT(n61971), .S0(buf_x[1232]), 
          .S1(buf_x[1233]));
    defparam add_4611_25.INIT0 = 16'h7888;
    defparam add_4611_25.INIT1 = 16'h7888;
    defparam add_4611_25.INJECT1_0 = "NO";
    defparam add_4611_25.INJECT1_1 = "NO";
    CCU2D add_4611_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[16]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[23]), .B1(nZ0_d2[16]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[17]), .CIN(n61969), .COUT(n61970), .S0(buf_x[1230]), 
          .S1(buf_x[1231]));
    defparam add_4611_23.INIT0 = 16'h7888;
    defparam add_4611_23.INIT1 = 16'h7888;
    defparam add_4611_23.INJECT1_0 = "NO";
    defparam add_4611_23.INJECT1_1 = "NO";
    CCU2D add_4611_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[16]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[21]), .B1(nZ0_d2[16]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[17]), .CIN(n61968), .COUT(n61969), .S0(buf_x[1228]), 
          .S1(buf_x[1229]));
    defparam add_4611_21.INIT0 = 16'h7888;
    defparam add_4611_21.INIT1 = 16'h7888;
    defparam add_4611_21.INJECT1_0 = "NO";
    defparam add_4611_21.INJECT1_1 = "NO";
    CCU2D add_4611_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[16]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[19]), .B1(nZ0_d2[16]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[17]), .CIN(n61967), .COUT(n61968), .S0(buf_x[1226]), 
          .S1(buf_x[1227]));
    defparam add_4611_19.INIT0 = 16'h7888;
    defparam add_4611_19.INIT1 = 16'h7888;
    defparam add_4611_19.INJECT1_0 = "NO";
    defparam add_4611_19.INJECT1_1 = "NO";
    CCU2D add_4611_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[16]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[17]), .B1(nZ0_d2[16]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[17]), .CIN(n61966), .COUT(n61967), .S0(buf_x[1224]), 
          .S1(buf_x[1225]));
    defparam add_4611_17.INIT0 = 16'h7888;
    defparam add_4611_17.INIT1 = 16'h7888;
    defparam add_4611_17.INJECT1_0 = "NO";
    defparam add_4611_17.INJECT1_1 = "NO";
    FD1S3AX buf_r_1299__500 (.D(buf_x[1299]), .CK(clock), .Q(buf_x[1650]));
    defparam buf_r_1299__500.GSR = "DISABLED";
    FD1S3AX buf_r_1298__501 (.D(buf_x[1298]), .CK(clock), .Q(buf_x[1649]));
    defparam buf_r_1298__501.GSR = "DISABLED";
    FD1S3AX buf_r_1297__502 (.D(buf_x[1297]), .CK(clock), .Q(buf_x[1648]));
    defparam buf_r_1297__502.GSR = "DISABLED";
    FD1S3AX buf_r_1296__503 (.D(buf_x[1296]), .CK(clock), .Q(buf_x[1647]));
    defparam buf_r_1296__503.GSR = "DISABLED";
    FD1S3AX buf_r_1295__504 (.D(buf_x[1295]), .CK(clock), .Q(buf_x[1646]));
    defparam buf_r_1295__504.GSR = "DISABLED";
    FD1S3AX buf_r_1294__505 (.D(buf_x[1294]), .CK(clock), .Q(buf_x[1645]));
    defparam buf_r_1294__505.GSR = "DISABLED";
    FD1S3AX buf_r_1293__506 (.D(buf_x[1293]), .CK(clock), .Q(buf_x[1644]));
    defparam buf_r_1293__506.GSR = "DISABLED";
    FD1S3AX buf_r_1292__507 (.D(buf_x[1292]), .CK(clock), .Q(buf_x[1643]));
    defparam buf_r_1292__507.GSR = "DISABLED";
    FD1S3AX buf_r_1291__508 (.D(buf_x[1291]), .CK(clock), .Q(buf_x[1642]));
    defparam buf_r_1291__508.GSR = "DISABLED";
    FD1S3AX buf_r_1290__509 (.D(buf_x[1290]), .CK(clock), .Q(buf_x[1641]));
    defparam buf_r_1290__509.GSR = "DISABLED";
    FD1S3AX buf_r_1289__510 (.D(buf_x[1289]), .CK(clock), .Q(buf_x[1640]));
    defparam buf_r_1289__510.GSR = "DISABLED";
    FD1S3AX buf_r_1288__511 (.D(buf_x[1288]), .CK(clock), .Q(buf_x[1639]));
    defparam buf_r_1288__511.GSR = "DISABLED";
    FD1S3AX buf_r_1287__512 (.D(buf_x[1287]), .CK(clock), .Q(buf_x[1638]));
    defparam buf_r_1287__512.GSR = "DISABLED";
    FD1S3AX buf_r_1286__513 (.D(buf_x[1286]), .CK(clock), .Q(buf_x[1637]));
    defparam buf_r_1286__513.GSR = "DISABLED";
    FD1S3AX buf_r_1285__514 (.D(buf_x[1285]), .CK(clock), .Q(buf_x[1636]));
    defparam buf_r_1285__514.GSR = "DISABLED";
    FD1S3AX buf_r_1284__515 (.D(buf_x[1284]), .CK(clock), .Q(buf_x[1635]));
    defparam buf_r_1284__515.GSR = "DISABLED";
    FD1S3AX buf_r_1283__516 (.D(buf_x[1283]), .CK(clock), .Q(buf_x[1634]));
    defparam buf_r_1283__516.GSR = "DISABLED";
    FD1S3AX buf_r_1282__517 (.D(buf_x[1282]), .CK(clock), .Q(buf_x[1633]));
    defparam buf_r_1282__517.GSR = "DISABLED";
    FD1S3AX buf_r_1281__518 (.D(buf_x[1281]), .CK(clock), .Q(buf_x[1632]));
    defparam buf_r_1281__518.GSR = "DISABLED";
    FD1S3AX buf_r_1280__519 (.D(buf_x[1280]), .CK(clock), .Q(buf_x[1631]));
    defparam buf_r_1280__519.GSR = "DISABLED";
    FD1S3AX buf_r_1279__520 (.D(buf_x[1279]), .CK(clock), .Q(buf_x[1630]));
    defparam buf_r_1279__520.GSR = "DISABLED";
    FD1S3AX buf_r_1278__521 (.D(buf_x[1278]), .CK(clock), .Q(buf_x[1629]));
    defparam buf_r_1278__521.GSR = "DISABLED";
    FD1S3AX buf_r_1277__522 (.D(buf_x[1277]), .CK(clock), .Q(buf_x[1628]));
    defparam buf_r_1277__522.GSR = "DISABLED";
    FD1S3AX buf_r_1276__523 (.D(buf_x[1276]), .CK(clock), .Q(buf_x[1627]));
    defparam buf_r_1276__523.GSR = "DISABLED";
    FD1S3AX buf_r_1275__524 (.D(buf_x[1275]), .CK(clock), .Q(buf_x[1626]));
    defparam buf_r_1275__524.GSR = "DISABLED";
    FD1S3AX buf_r_1274__525 (.D(buf_x[1274]), .CK(clock), .Q(buf_x[1625]));
    defparam buf_r_1274__525.GSR = "DISABLED";
    FD1S3AX buf_r_1273__526 (.D(buf_x[1273]), .CK(clock), .Q(buf_x[1624]));
    defparam buf_r_1273__526.GSR = "DISABLED";
    FD1S3AX buf_r_1272__527 (.D(buf_x[1272]), .CK(clock), .Q(buf_x[1623]));
    defparam buf_r_1272__527.GSR = "DISABLED";
    FD1S3AX buf_r_1271__528 (.D(buf_x[1271]), .CK(clock), .Q(buf_x[1622]));
    defparam buf_r_1271__528.GSR = "DISABLED";
    FD1S3AX buf_r_1268__531 (.D(buf_x[1268]), .CK(clock), .Q(buf_r[1268]));
    defparam buf_r_1268__531.GSR = "DISABLED";
    FD1S3AX buf_r_1267__532 (.D(buf_x[1267]), .CK(clock), .Q(buf_r[1267]));
    defparam buf_r_1267__532.GSR = "DISABLED";
    FD1S3AX buf_r_1266__533 (.D(buf_x[1266]), .CK(clock), .Q(buf_r[1266]));
    defparam buf_r_1266__533.GSR = "DISABLED";
    FD1S3AX buf_r_1265__534 (.D(buf_x[1265]), .CK(clock), .Q(buf_r[1265]));
    defparam buf_r_1265__534.GSR = "DISABLED";
    FD1S3AX buf_r_1264__535 (.D(buf_x[1264]), .CK(clock), .Q(buf_r[1264]));
    defparam buf_r_1264__535.GSR = "DISABLED";
    FD1S3AX buf_r_1263__536 (.D(buf_x[1263]), .CK(clock), .Q(buf_r[1263]));
    defparam buf_r_1263__536.GSR = "DISABLED";
    FD1S3AX buf_r_1262__537 (.D(buf_x[1262]), .CK(clock), .Q(buf_r[1262]));
    defparam buf_r_1262__537.GSR = "DISABLED";
    FD1S3AX buf_r_1261__538 (.D(buf_x[1261]), .CK(clock), .Q(buf_r[1261]));
    defparam buf_r_1261__538.GSR = "DISABLED";
    FD1S3AX buf_r_1260__539 (.D(buf_x[1260]), .CK(clock), .Q(buf_r[1260]));
    defparam buf_r_1260__539.GSR = "DISABLED";
    FD1S3AX buf_r_1259__540 (.D(buf_x[1259]), .CK(clock), .Q(buf_r[1259]));
    defparam buf_r_1259__540.GSR = "DISABLED";
    FD1S3AX buf_r_1258__541 (.D(buf_x[1258]), .CK(clock), .Q(buf_r[1258]));
    defparam buf_r_1258__541.GSR = "DISABLED";
    FD1S3AX buf_r_1257__542 (.D(buf_x[1257]), .CK(clock), .Q(buf_r[1257]));
    defparam buf_r_1257__542.GSR = "DISABLED";
    FD1S3AX buf_r_1256__543 (.D(buf_x[1256]), .CK(clock), .Q(buf_r[1256]));
    defparam buf_r_1256__543.GSR = "DISABLED";
    FD1S3AX buf_r_1255__544 (.D(buf_x[1255]), .CK(clock), .Q(buf_r[1255]));
    defparam buf_r_1255__544.GSR = "DISABLED";
    FD1S3AX buf_r_1254__545 (.D(buf_x[1254]), .CK(clock), .Q(buf_r[1254]));
    defparam buf_r_1254__545.GSR = "DISABLED";
    FD1S3AX buf_r_1253__546 (.D(buf_x[1253]), .CK(clock), .Q(buf_r[1253]));
    defparam buf_r_1253__546.GSR = "DISABLED";
    FD1S3AX buf_r_1252__547 (.D(buf_x[1252]), .CK(clock), .Q(buf_r[1252]));
    defparam buf_r_1252__547.GSR = "DISABLED";
    FD1S3AX buf_r_1251__548 (.D(buf_x[1251]), .CK(clock), .Q(buf_r[1251]));
    defparam buf_r_1251__548.GSR = "DISABLED";
    FD1S3AX buf_r_1250__549 (.D(buf_x[1250]), .CK(clock), .Q(buf_r[1250]));
    defparam buf_r_1250__549.GSR = "DISABLED";
    FD1S3AX buf_r_1249__550 (.D(buf_x[1249]), .CK(clock), .Q(buf_r[1249]));
    defparam buf_r_1249__550.GSR = "DISABLED";
    FD1S3AX buf_r_1248__551 (.D(buf_x[1248]), .CK(clock), .Q(buf_r[1248]));
    defparam buf_r_1248__551.GSR = "DISABLED";
    FD1S3AX buf_r_1247__552 (.D(buf_x[1247]), .CK(clock), .Q(buf_r[1247]));
    defparam buf_r_1247__552.GSR = "DISABLED";
    FD1S3AX buf_r_1246__553 (.D(buf_x[1246]), .CK(clock), .Q(buf_r[1246]));
    defparam buf_r_1246__553.GSR = "DISABLED";
    FD1S3AX buf_r_1245__554 (.D(buf_x[1245]), .CK(clock), .Q(buf_r[1245]));
    defparam buf_r_1245__554.GSR = "DISABLED";
    FD1S3AX buf_r_1244__555 (.D(buf_x[1244]), .CK(clock), .Q(buf_r[1244]));
    defparam buf_r_1244__555.GSR = "DISABLED";
    FD1S3AX buf_r_1243__556 (.D(buf_x[1243]), .CK(clock), .Q(buf_r[1243]));
    defparam buf_r_1243__556.GSR = "DISABLED";
    FD1S3AX buf_r_1242__557 (.D(buf_x[1242]), .CK(clock), .Q(buf_r[1242]));
    defparam buf_r_1242__557.GSR = "DISABLED";
    FD1S3AX buf_r_1241__558 (.D(buf_x[1241]), .CK(clock), .Q(buf_r[1241]));
    defparam buf_r_1241__558.GSR = "DISABLED";
    FD1S3AX buf_r_1240__559 (.D(buf_x[1240]), .CK(clock), .Q(buf_r[1240]));
    defparam buf_r_1240__559.GSR = "DISABLED";
    FD1S3AX buf_r_1237__562 (.D(buf_x[1237]), .CK(clock), .Q(buf_r[1237]));
    defparam buf_r_1237__562.GSR = "DISABLED";
    FD1S3AX buf_r_1236__563 (.D(buf_x[1236]), .CK(clock), .Q(buf_r[1236]));
    defparam buf_r_1236__563.GSR = "DISABLED";
    FD1S3AX buf_r_1235__564 (.D(buf_x[1235]), .CK(clock), .Q(buf_r[1235]));
    defparam buf_r_1235__564.GSR = "DISABLED";
    FD1S3AX buf_r_1234__565 (.D(buf_x[1234]), .CK(clock), .Q(buf_r[1234]));
    defparam buf_r_1234__565.GSR = "DISABLED";
    FD1S3AX buf_r_1233__566 (.D(buf_x[1233]), .CK(clock), .Q(buf_r[1233]));
    defparam buf_r_1233__566.GSR = "DISABLED";
    FD1S3AX buf_r_1232__567 (.D(buf_x[1232]), .CK(clock), .Q(buf_r[1232]));
    defparam buf_r_1232__567.GSR = "DISABLED";
    FD1S3AX buf_r_1231__568 (.D(buf_x[1231]), .CK(clock), .Q(buf_r[1231]));
    defparam buf_r_1231__568.GSR = "DISABLED";
    FD1S3AX buf_r_1230__569 (.D(buf_x[1230]), .CK(clock), .Q(buf_r[1230]));
    defparam buf_r_1230__569.GSR = "DISABLED";
    FD1S3AX buf_r_1229__570 (.D(buf_x[1229]), .CK(clock), .Q(buf_r[1229]));
    defparam buf_r_1229__570.GSR = "DISABLED";
    FD1S3AX buf_r_1228__571 (.D(buf_x[1228]), .CK(clock), .Q(buf_r[1228]));
    defparam buf_r_1228__571.GSR = "DISABLED";
    FD1S3AX buf_r_1227__572 (.D(buf_x[1227]), .CK(clock), .Q(buf_r[1227]));
    defparam buf_r_1227__572.GSR = "DISABLED";
    FD1S3AX buf_r_1226__573 (.D(buf_x[1226]), .CK(clock), .Q(buf_r[1226]));
    defparam buf_r_1226__573.GSR = "DISABLED";
    FD1S3AX buf_r_1225__574 (.D(buf_x[1225]), .CK(clock), .Q(buf_r[1225]));
    defparam buf_r_1225__574.GSR = "DISABLED";
    FD1S3AX buf_r_1224__575 (.D(buf_x[1224]), .CK(clock), .Q(buf_r[1224]));
    defparam buf_r_1224__575.GSR = "DISABLED";
    FD1S3AX buf_r_1223__576 (.D(buf_x[1223]), .CK(clock), .Q(buf_r[1223]));
    defparam buf_r_1223__576.GSR = "DISABLED";
    FD1S3AX buf_r_1222__577 (.D(buf_x[1222]), .CK(clock), .Q(buf_r[1222]));
    defparam buf_r_1222__577.GSR = "DISABLED";
    FD1S3AX buf_r_1221__578 (.D(buf_x[1221]), .CK(clock), .Q(buf_r[1221]));
    defparam buf_r_1221__578.GSR = "DISABLED";
    FD1S3AX buf_r_1220__579 (.D(buf_x[1220]), .CK(clock), .Q(buf_r[1220]));
    defparam buf_r_1220__579.GSR = "DISABLED";
    FD1S3AX buf_r_1219__580 (.D(buf_x[1219]), .CK(clock), .Q(buf_r[1219]));
    defparam buf_r_1219__580.GSR = "DISABLED";
    FD1S3AX buf_r_1218__581 (.D(buf_x[1218]), .CK(clock), .Q(buf_r[1218]));
    defparam buf_r_1218__581.GSR = "DISABLED";
    FD1S3AX buf_r_1217__582 (.D(buf_x[1217]), .CK(clock), .Q(buf_r[1217]));
    defparam buf_r_1217__582.GSR = "DISABLED";
    FD1S3AX buf_r_1216__583 (.D(buf_x[1216]), .CK(clock), .Q(buf_r[1216]));
    defparam buf_r_1216__583.GSR = "DISABLED";
    FD1S3AX buf_r_1215__584 (.D(buf_x[1215]), .CK(clock), .Q(buf_r[1215]));
    defparam buf_r_1215__584.GSR = "DISABLED";
    FD1S3AX buf_r_1214__585 (.D(buf_x[1214]), .CK(clock), .Q(buf_r[1214]));
    defparam buf_r_1214__585.GSR = "DISABLED";
    FD1S3AX buf_r_1213__586 (.D(buf_x[1213]), .CK(clock), .Q(buf_r[1213]));
    defparam buf_r_1213__586.GSR = "DISABLED";
    FD1S3AX buf_r_1212__587 (.D(buf_x[1212]), .CK(clock), .Q(buf_r[1212]));
    defparam buf_r_1212__587.GSR = "DISABLED";
    FD1S3AX buf_r_1211__588 (.D(buf_x[1211]), .CK(clock), .Q(buf_r[1211]));
    defparam buf_r_1211__588.GSR = "DISABLED";
    FD1S3AX buf_r_1210__589 (.D(buf_x[1210]), .CK(clock), .Q(buf_r[1210]));
    defparam buf_r_1210__589.GSR = "DISABLED";
    FD1S3AX buf_r_1209__590 (.D(buf_x[1209]), .CK(clock), .Q(buf_x[1795]));
    defparam buf_r_1209__590.GSR = "DISABLED";
    FD1S3AX buf_r_1206__593 (.D(buf_x[1206]), .CK(clock), .Q(buf_r[1206]));
    defparam buf_r_1206__593.GSR = "DISABLED";
    FD1S3AX buf_r_1205__594 (.D(buf_x[1205]), .CK(clock), .Q(buf_r[1205]));
    defparam buf_r_1205__594.GSR = "DISABLED";
    FD1S3AX buf_r_1204__595 (.D(buf_x[1204]), .CK(clock), .Q(buf_r[1204]));
    defparam buf_r_1204__595.GSR = "DISABLED";
    FD1S3AX buf_r_1203__596 (.D(buf_x[1203]), .CK(clock), .Q(buf_r[1203]));
    defparam buf_r_1203__596.GSR = "DISABLED";
    FD1S3AX buf_r_1202__597 (.D(buf_x[1202]), .CK(clock), .Q(buf_r[1202]));
    defparam buf_r_1202__597.GSR = "DISABLED";
    FD1S3AX buf_r_1201__598 (.D(buf_x[1201]), .CK(clock), .Q(buf_r[1201]));
    defparam buf_r_1201__598.GSR = "DISABLED";
    FD1S3AX buf_r_1200__599 (.D(buf_x[1200]), .CK(clock), .Q(buf_r[1200]));
    defparam buf_r_1200__599.GSR = "DISABLED";
    FD1S3AX buf_r_1199__600 (.D(buf_x[1199]), .CK(clock), .Q(buf_r[1199]));
    defparam buf_r_1199__600.GSR = "DISABLED";
    FD1S3AX buf_r_1198__601 (.D(buf_x[1198]), .CK(clock), .Q(buf_r[1198]));
    defparam buf_r_1198__601.GSR = "DISABLED";
    FD1S3AX buf_r_1197__602 (.D(buf_x[1197]), .CK(clock), .Q(buf_r[1197]));
    defparam buf_r_1197__602.GSR = "DISABLED";
    FD1S3AX buf_r_1196__603 (.D(buf_x[1196]), .CK(clock), .Q(buf_r[1196]));
    defparam buf_r_1196__603.GSR = "DISABLED";
    FD1S3AX buf_r_1195__604 (.D(buf_x[1195]), .CK(clock), .Q(buf_r[1195]));
    defparam buf_r_1195__604.GSR = "DISABLED";
    FD1S3AX buf_r_1194__605 (.D(buf_x[1194]), .CK(clock), .Q(buf_r[1194]));
    defparam buf_r_1194__605.GSR = "DISABLED";
    FD1S3AX buf_r_1193__606 (.D(buf_x[1193]), .CK(clock), .Q(buf_r[1193]));
    defparam buf_r_1193__606.GSR = "DISABLED";
    FD1S3AX buf_r_1192__607 (.D(buf_x[1192]), .CK(clock), .Q(buf_r[1192]));
    defparam buf_r_1192__607.GSR = "DISABLED";
    FD1S3AX buf_r_1191__608 (.D(buf_x[1191]), .CK(clock), .Q(buf_r[1191]));
    defparam buf_r_1191__608.GSR = "DISABLED";
    FD1S3AX buf_r_1190__609 (.D(buf_x[1190]), .CK(clock), .Q(buf_r[1190]));
    defparam buf_r_1190__609.GSR = "DISABLED";
    FD1S3AX buf_r_1189__610 (.D(buf_x[1189]), .CK(clock), .Q(buf_r[1189]));
    defparam buf_r_1189__610.GSR = "DISABLED";
    FD1S3AX buf_r_1188__611 (.D(buf_x[1188]), .CK(clock), .Q(buf_r[1188]));
    defparam buf_r_1188__611.GSR = "DISABLED";
    FD1S3AX buf_r_1187__612 (.D(buf_x[1187]), .CK(clock), .Q(buf_r[1187]));
    defparam buf_r_1187__612.GSR = "DISABLED";
    FD1S3AX buf_r_1186__613 (.D(buf_x[1186]), .CK(clock), .Q(buf_r[1186]));
    defparam buf_r_1186__613.GSR = "DISABLED";
    FD1S3AX buf_r_1185__614 (.D(buf_x[1185]), .CK(clock), .Q(buf_r[1185]));
    defparam buf_r_1185__614.GSR = "DISABLED";
    FD1S3AX buf_r_1184__615 (.D(buf_x[1184]), .CK(clock), .Q(buf_r[1184]));
    defparam buf_r_1184__615.GSR = "DISABLED";
    FD1S3AX buf_r_1183__616 (.D(buf_x[1183]), .CK(clock), .Q(buf_r[1183]));
    defparam buf_r_1183__616.GSR = "DISABLED";
    FD1S3AX buf_r_1182__617 (.D(buf_x[1182]), .CK(clock), .Q(buf_r[1182]));
    defparam buf_r_1182__617.GSR = "DISABLED";
    FD1S3AX buf_r_1181__618 (.D(buf_x[1181]), .CK(clock), .Q(buf_r[1181]));
    defparam buf_r_1181__618.GSR = "DISABLED";
    FD1S3AX buf_r_1180__619 (.D(buf_x[1180]), .CK(clock), .Q(buf_r[1180]));
    defparam buf_r_1180__619.GSR = "DISABLED";
    FD1S3AX buf_r_1179__620 (.D(buf_x[1179]), .CK(clock), .Q(buf_r[1179]));
    defparam buf_r_1179__620.GSR = "DISABLED";
    FD1S3AX buf_r_1178__621 (.D(buf_x[1178]), .CK(clock), .Q(buf_r[1178]));
    defparam buf_r_1178__621.GSR = "DISABLED";
    FD1S3AX buf_r_1175__624 (.D(buf_x[1175]), .CK(clock), .Q(buf_r[1175]));
    defparam buf_r_1175__624.GSR = "DISABLED";
    FD1S3AX buf_r_1174__625 (.D(buf_x[1174]), .CK(clock), .Q(buf_r[1174]));
    defparam buf_r_1174__625.GSR = "DISABLED";
    FD1S3AX buf_r_1173__626 (.D(buf_x[1173]), .CK(clock), .Q(buf_r[1173]));
    defparam buf_r_1173__626.GSR = "DISABLED";
    FD1S3AX buf_r_1172__627 (.D(buf_x[1172]), .CK(clock), .Q(buf_r[1172]));
    defparam buf_r_1172__627.GSR = "DISABLED";
    FD1S3AX buf_r_1171__628 (.D(buf_x[1171]), .CK(clock), .Q(buf_r[1171]));
    defparam buf_r_1171__628.GSR = "DISABLED";
    FD1S3AX buf_r_1170__629 (.D(buf_x[1170]), .CK(clock), .Q(buf_r[1170]));
    defparam buf_r_1170__629.GSR = "DISABLED";
    FD1S3AX buf_r_1169__630 (.D(buf_x[1169]), .CK(clock), .Q(buf_r[1169]));
    defparam buf_r_1169__630.GSR = "DISABLED";
    FD1S3AX buf_r_1168__631 (.D(buf_x[1168]), .CK(clock), .Q(buf_r[1168]));
    defparam buf_r_1168__631.GSR = "DISABLED";
    FD1S3AX buf_r_1167__632 (.D(buf_x[1167]), .CK(clock), .Q(buf_r[1167]));
    defparam buf_r_1167__632.GSR = "DISABLED";
    FD1S3AX buf_r_1166__633 (.D(buf_x[1166]), .CK(clock), .Q(buf_r[1166]));
    defparam buf_r_1166__633.GSR = "DISABLED";
    FD1S3AX buf_r_1165__634 (.D(buf_x[1165]), .CK(clock), .Q(buf_r[1165]));
    defparam buf_r_1165__634.GSR = "DISABLED";
    FD1S3AX buf_r_1164__635 (.D(buf_x[1164]), .CK(clock), .Q(buf_r[1164]));
    defparam buf_r_1164__635.GSR = "DISABLED";
    FD1S3AX buf_r_1163__636 (.D(buf_x[1163]), .CK(clock), .Q(buf_r[1163]));
    defparam buf_r_1163__636.GSR = "DISABLED";
    FD1S3AX buf_r_1162__637 (.D(buf_x[1162]), .CK(clock), .Q(buf_r[1162]));
    defparam buf_r_1162__637.GSR = "DISABLED";
    FD1S3AX buf_r_1161__638 (.D(buf_x[1161]), .CK(clock), .Q(buf_r[1161]));
    defparam buf_r_1161__638.GSR = "DISABLED";
    FD1S3AX buf_r_1160__639 (.D(buf_x[1160]), .CK(clock), .Q(buf_r[1160]));
    defparam buf_r_1160__639.GSR = "DISABLED";
    FD1S3AX buf_r_1159__640 (.D(buf_x[1159]), .CK(clock), .Q(buf_r[1159]));
    defparam buf_r_1159__640.GSR = "DISABLED";
    FD1S3AX buf_r_1158__641 (.D(buf_x[1158]), .CK(clock), .Q(buf_r[1158]));
    defparam buf_r_1158__641.GSR = "DISABLED";
    FD1S3AX buf_r_1157__642 (.D(buf_x[1157]), .CK(clock), .Q(buf_r[1157]));
    defparam buf_r_1157__642.GSR = "DISABLED";
    FD1S3AX buf_r_1156__643 (.D(buf_x[1156]), .CK(clock), .Q(buf_r[1156]));
    defparam buf_r_1156__643.GSR = "DISABLED";
    FD1S3AX buf_r_1155__644 (.D(buf_x[1155]), .CK(clock), .Q(buf_r[1155]));
    defparam buf_r_1155__644.GSR = "DISABLED";
    FD1S3AX buf_r_1154__645 (.D(buf_x[1154]), .CK(clock), .Q(buf_r[1154]));
    defparam buf_r_1154__645.GSR = "DISABLED";
    FD1S3AX buf_r_1153__646 (.D(buf_x[1153]), .CK(clock), .Q(buf_r[1153]));
    defparam buf_r_1153__646.GSR = "DISABLED";
    FD1S3AX buf_r_1152__647 (.D(buf_x[1152]), .CK(clock), .Q(buf_r[1152]));
    defparam buf_r_1152__647.GSR = "DISABLED";
    FD1S3AX buf_r_1151__648 (.D(buf_x[1151]), .CK(clock), .Q(buf_r[1151]));
    defparam buf_r_1151__648.GSR = "DISABLED";
    FD1S3AX buf_r_1150__649 (.D(buf_x[1150]), .CK(clock), .Q(buf_r[1150]));
    defparam buf_r_1150__649.GSR = "DISABLED";
    FD1S3AX buf_r_1149__650 (.D(buf_x[1149]), .CK(clock), .Q(buf_r[1149]));
    defparam buf_r_1149__650.GSR = "DISABLED";
    FD1S3AX buf_r_1148__651 (.D(buf_x[1148]), .CK(clock), .Q(buf_r[1148]));
    defparam buf_r_1148__651.GSR = "DISABLED";
    FD1S3AX buf_r_1147__652 (.D(buf_x[1147]), .CK(clock), .Q(buf_x[1556]));
    defparam buf_r_1147__652.GSR = "DISABLED";
    FD1S3AX buf_r_1144__655 (.D(buf_x[1144]), .CK(clock), .Q(buf_r[1144]));
    defparam buf_r_1144__655.GSR = "DISABLED";
    FD1S3AX buf_r_1143__656 (.D(buf_x[1143]), .CK(clock), .Q(buf_r[1143]));
    defparam buf_r_1143__656.GSR = "DISABLED";
    FD1S3AX buf_r_1142__657 (.D(buf_x[1142]), .CK(clock), .Q(buf_r[1142]));
    defparam buf_r_1142__657.GSR = "DISABLED";
    FD1S3AX buf_r_1141__658 (.D(buf_x[1141]), .CK(clock), .Q(buf_r[1141]));
    defparam buf_r_1141__658.GSR = "DISABLED";
    FD1S3AX buf_r_1140__659 (.D(buf_x[1140]), .CK(clock), .Q(buf_r[1140]));
    defparam buf_r_1140__659.GSR = "DISABLED";
    FD1S3AX buf_r_1139__660 (.D(buf_x[1139]), .CK(clock), .Q(buf_r[1139]));
    defparam buf_r_1139__660.GSR = "DISABLED";
    FD1S3AX buf_r_1138__661 (.D(buf_x[1138]), .CK(clock), .Q(buf_r[1138]));
    defparam buf_r_1138__661.GSR = "DISABLED";
    FD1S3AX buf_r_1137__662 (.D(buf_x[1137]), .CK(clock), .Q(buf_r[1137]));
    defparam buf_r_1137__662.GSR = "DISABLED";
    FD1S3AX buf_r_1136__663 (.D(buf_x[1136]), .CK(clock), .Q(buf_r[1136]));
    defparam buf_r_1136__663.GSR = "DISABLED";
    FD1S3AX buf_r_1135__664 (.D(buf_x[1135]), .CK(clock), .Q(buf_r[1135]));
    defparam buf_r_1135__664.GSR = "DISABLED";
    FD1S3AX buf_r_1134__665 (.D(buf_x[1134]), .CK(clock), .Q(buf_r[1134]));
    defparam buf_r_1134__665.GSR = "DISABLED";
    FD1S3AX buf_r_1133__666 (.D(buf_x[1133]), .CK(clock), .Q(buf_r[1133]));
    defparam buf_r_1133__666.GSR = "DISABLED";
    FD1S3AX buf_r_1132__667 (.D(buf_x[1132]), .CK(clock), .Q(buf_r[1132]));
    defparam buf_r_1132__667.GSR = "DISABLED";
    FD1S3AX buf_r_1131__668 (.D(buf_x[1131]), .CK(clock), .Q(buf_r[1131]));
    defparam buf_r_1131__668.GSR = "DISABLED";
    FD1S3AX buf_r_1130__669 (.D(buf_x[1130]), .CK(clock), .Q(buf_r[1130]));
    defparam buf_r_1130__669.GSR = "DISABLED";
    FD1S3AX buf_r_1129__670 (.D(buf_x[1129]), .CK(clock), .Q(buf_r[1129]));
    defparam buf_r_1129__670.GSR = "DISABLED";
    FD1S3AX buf_r_1128__671 (.D(buf_x[1128]), .CK(clock), .Q(buf_r[1128]));
    defparam buf_r_1128__671.GSR = "DISABLED";
    FD1S3AX buf_r_1127__672 (.D(buf_x[1127]), .CK(clock), .Q(buf_r[1127]));
    defparam buf_r_1127__672.GSR = "DISABLED";
    FD1S3AX buf_r_1126__673 (.D(buf_x[1126]), .CK(clock), .Q(buf_r[1126]));
    defparam buf_r_1126__673.GSR = "DISABLED";
    FD1S3AX buf_r_1125__674 (.D(buf_x[1125]), .CK(clock), .Q(buf_r[1125]));
    defparam buf_r_1125__674.GSR = "DISABLED";
    FD1S3AX buf_r_1124__675 (.D(buf_x[1124]), .CK(clock), .Q(buf_r[1124]));
    defparam buf_r_1124__675.GSR = "DISABLED";
    FD1S3AX buf_r_1123__676 (.D(buf_x[1123]), .CK(clock), .Q(buf_r[1123]));
    defparam buf_r_1123__676.GSR = "DISABLED";
    FD1S3AX buf_r_1122__677 (.D(buf_x[1122]), .CK(clock), .Q(buf_r[1122]));
    defparam buf_r_1122__677.GSR = "DISABLED";
    FD1S3AX buf_r_1121__678 (.D(buf_x[1121]), .CK(clock), .Q(buf_r[1121]));
    defparam buf_r_1121__678.GSR = "DISABLED";
    FD1S3AX buf_r_1120__679 (.D(buf_x[1120]), .CK(clock), .Q(buf_r[1120]));
    defparam buf_r_1120__679.GSR = "DISABLED";
    FD1S3AX buf_r_1119__680 (.D(buf_x[1119]), .CK(clock), .Q(buf_r[1119]));
    defparam buf_r_1119__680.GSR = "DISABLED";
    FD1S3AX buf_r_1118__681 (.D(buf_x[1118]), .CK(clock), .Q(buf_r[1118]));
    defparam buf_r_1118__681.GSR = "DISABLED";
    FD1S3AX buf_r_1117__682 (.D(buf_x[1117]), .CK(clock), .Q(buf_r[1117]));
    defparam buf_r_1117__682.GSR = "DISABLED";
    FD1S3AX buf_r_1116__683 (.D(buf_x[1116]), .CK(clock), .Q(buf_r[1116]));
    defparam buf_r_1116__683.GSR = "DISABLED";
    FD1S3AX buf_r_1113__686 (.D(buf_x[1113]), .CK(clock), .Q(buf_r[1113]));
    defparam buf_r_1113__686.GSR = "DISABLED";
    FD1S3AX buf_r_1112__687 (.D(buf_x[1112]), .CK(clock), .Q(buf_r[1112]));
    defparam buf_r_1112__687.GSR = "DISABLED";
    FD1S3AX buf_r_1111__688 (.D(buf_x[1111]), .CK(clock), .Q(buf_r[1111]));
    defparam buf_r_1111__688.GSR = "DISABLED";
    FD1S3AX buf_r_1110__689 (.D(buf_x[1110]), .CK(clock), .Q(buf_r[1110]));
    defparam buf_r_1110__689.GSR = "DISABLED";
    FD1S3AX buf_r_1109__690 (.D(buf_x[1109]), .CK(clock), .Q(buf_r[1109]));
    defparam buf_r_1109__690.GSR = "DISABLED";
    FD1S3AX buf_r_1108__691 (.D(buf_x[1108]), .CK(clock), .Q(buf_r[1108]));
    defparam buf_r_1108__691.GSR = "DISABLED";
    FD1S3AX buf_r_1107__692 (.D(buf_x[1107]), .CK(clock), .Q(buf_r[1107]));
    defparam buf_r_1107__692.GSR = "DISABLED";
    FD1S3AX buf_r_1106__693 (.D(buf_x[1106]), .CK(clock), .Q(buf_r[1106]));
    defparam buf_r_1106__693.GSR = "DISABLED";
    FD1S3AX buf_r_1105__694 (.D(buf_x[1105]), .CK(clock), .Q(buf_r[1105]));
    defparam buf_r_1105__694.GSR = "DISABLED";
    FD1S3AX buf_r_1104__695 (.D(buf_x[1104]), .CK(clock), .Q(buf_r[1104]));
    defparam buf_r_1104__695.GSR = "DISABLED";
    FD1S3AX buf_r_1103__696 (.D(buf_x[1103]), .CK(clock), .Q(buf_r[1103]));
    defparam buf_r_1103__696.GSR = "DISABLED";
    FD1S3AX buf_r_1102__697 (.D(buf_x[1102]), .CK(clock), .Q(buf_r[1102]));
    defparam buf_r_1102__697.GSR = "DISABLED";
    FD1S3AX buf_r_1101__698 (.D(buf_x[1101]), .CK(clock), .Q(buf_r[1101]));
    defparam buf_r_1101__698.GSR = "DISABLED";
    FD1S3AX buf_r_1100__699 (.D(buf_x[1100]), .CK(clock), .Q(buf_r[1100]));
    defparam buf_r_1100__699.GSR = "DISABLED";
    FD1S3AX buf_r_1099__700 (.D(buf_x[1099]), .CK(clock), .Q(buf_r[1099]));
    defparam buf_r_1099__700.GSR = "DISABLED";
    FD1S3AX buf_r_1098__701 (.D(buf_x[1098]), .CK(clock), .Q(buf_r[1098]));
    defparam buf_r_1098__701.GSR = "DISABLED";
    FD1S3AX buf_r_1097__702 (.D(buf_x[1097]), .CK(clock), .Q(buf_r[1097]));
    defparam buf_r_1097__702.GSR = "DISABLED";
    FD1S3AX buf_r_1096__703 (.D(buf_x[1096]), .CK(clock), .Q(buf_r[1096]));
    defparam buf_r_1096__703.GSR = "DISABLED";
    FD1S3AX buf_r_1095__704 (.D(buf_x[1095]), .CK(clock), .Q(buf_r[1095]));
    defparam buf_r_1095__704.GSR = "DISABLED";
    FD1S3AX buf_r_1094__705 (.D(buf_x[1094]), .CK(clock), .Q(buf_r[1094]));
    defparam buf_r_1094__705.GSR = "DISABLED";
    FD1S3AX buf_r_1093__706 (.D(buf_x[1093]), .CK(clock), .Q(buf_r[1093]));
    defparam buf_r_1093__706.GSR = "DISABLED";
    FD1S3AX buf_r_1092__707 (.D(buf_x[1092]), .CK(clock), .Q(buf_r[1092]));
    defparam buf_r_1092__707.GSR = "DISABLED";
    FD1S3AX buf_r_1091__708 (.D(buf_x[1091]), .CK(clock), .Q(buf_r[1091]));
    defparam buf_r_1091__708.GSR = "DISABLED";
    FD1S3AX buf_r_1090__709 (.D(buf_x[1090]), .CK(clock), .Q(buf_r[1090]));
    defparam buf_r_1090__709.GSR = "DISABLED";
    FD1S3AX buf_r_1089__710 (.D(buf_x[1089]), .CK(clock), .Q(buf_r[1089]));
    defparam buf_r_1089__710.GSR = "DISABLED";
    FD1S3AX buf_r_1088__711 (.D(buf_x[1088]), .CK(clock), .Q(buf_r[1088]));
    defparam buf_r_1088__711.GSR = "DISABLED";
    FD1S3AX buf_r_1087__712 (.D(buf_x[1087]), .CK(clock), .Q(buf_r[1087]));
    defparam buf_r_1087__712.GSR = "DISABLED";
    FD1S3AX buf_r_1086__713 (.D(buf_x[1086]), .CK(clock), .Q(buf_r[1086]));
    defparam buf_r_1086__713.GSR = "DISABLED";
    FD1S3AX buf_r_1085__714 (.D(buf_x[1085]), .CK(clock), .Q(buf_x[1758]));
    defparam buf_r_1085__714.GSR = "DISABLED";
    FD1S3AX buf_r_1082__717 (.D(buf_x[1082]), .CK(clock), .Q(buf_r[1082]));
    defparam buf_r_1082__717.GSR = "DISABLED";
    FD1S3AX buf_r_1081__718 (.D(buf_x[1081]), .CK(clock), .Q(buf_r[1081]));
    defparam buf_r_1081__718.GSR = "DISABLED";
    FD1S3AX buf_r_1080__719 (.D(buf_x[1080]), .CK(clock), .Q(buf_r[1080]));
    defparam buf_r_1080__719.GSR = "DISABLED";
    FD1S3AX buf_r_1079__720 (.D(buf_x[1079]), .CK(clock), .Q(buf_r[1079]));
    defparam buf_r_1079__720.GSR = "DISABLED";
    FD1S3AX buf_r_1078__721 (.D(buf_x[1078]), .CK(clock), .Q(buf_r[1078]));
    defparam buf_r_1078__721.GSR = "DISABLED";
    FD1S3AX buf_r_1077__722 (.D(buf_x[1077]), .CK(clock), .Q(buf_r[1077]));
    defparam buf_r_1077__722.GSR = "DISABLED";
    FD1S3AX buf_r_1076__723 (.D(buf_x[1076]), .CK(clock), .Q(buf_r[1076]));
    defparam buf_r_1076__723.GSR = "DISABLED";
    FD1S3AX buf_r_1075__724 (.D(buf_x[1075]), .CK(clock), .Q(buf_r[1075]));
    defparam buf_r_1075__724.GSR = "DISABLED";
    FD1S3AX buf_r_1074__725 (.D(buf_x[1074]), .CK(clock), .Q(buf_r[1074]));
    defparam buf_r_1074__725.GSR = "DISABLED";
    FD1S3AX buf_r_1073__726 (.D(buf_x[1073]), .CK(clock), .Q(buf_r[1073]));
    defparam buf_r_1073__726.GSR = "DISABLED";
    FD1S3AX buf_r_1072__727 (.D(buf_x[1072]), .CK(clock), .Q(buf_r[1072]));
    defparam buf_r_1072__727.GSR = "DISABLED";
    FD1S3AX buf_r_1071__728 (.D(buf_x[1071]), .CK(clock), .Q(buf_r[1071]));
    defparam buf_r_1071__728.GSR = "DISABLED";
    FD1S3AX buf_r_1070__729 (.D(buf_x[1070]), .CK(clock), .Q(buf_r[1070]));
    defparam buf_r_1070__729.GSR = "DISABLED";
    FD1S3AX buf_r_1069__730 (.D(buf_x[1069]), .CK(clock), .Q(buf_r[1069]));
    defparam buf_r_1069__730.GSR = "DISABLED";
    FD1S3AX buf_r_1068__731 (.D(buf_x[1068]), .CK(clock), .Q(buf_r[1068]));
    defparam buf_r_1068__731.GSR = "DISABLED";
    FD1S3AX buf_r_1067__732 (.D(buf_x[1067]), .CK(clock), .Q(buf_r[1067]));
    defparam buf_r_1067__732.GSR = "DISABLED";
    FD1S3AX buf_r_1066__733 (.D(buf_x[1066]), .CK(clock), .Q(buf_r[1066]));
    defparam buf_r_1066__733.GSR = "DISABLED";
    FD1S3AX buf_r_1065__734 (.D(buf_x[1065]), .CK(clock), .Q(buf_r[1065]));
    defparam buf_r_1065__734.GSR = "DISABLED";
    FD1S3AX buf_r_1064__735 (.D(buf_x[1064]), .CK(clock), .Q(buf_r[1064]));
    defparam buf_r_1064__735.GSR = "DISABLED";
    FD1S3AX buf_r_1063__736 (.D(buf_x[1063]), .CK(clock), .Q(buf_r[1063]));
    defparam buf_r_1063__736.GSR = "DISABLED";
    FD1S3AX buf_r_1062__737 (.D(buf_x[1062]), .CK(clock), .Q(buf_r[1062]));
    defparam buf_r_1062__737.GSR = "DISABLED";
    FD1S3AX buf_r_1061__738 (.D(buf_x[1061]), .CK(clock), .Q(buf_r[1061]));
    defparam buf_r_1061__738.GSR = "DISABLED";
    FD1S3AX buf_r_1060__739 (.D(buf_x[1060]), .CK(clock), .Q(buf_r[1060]));
    defparam buf_r_1060__739.GSR = "DISABLED";
    FD1S3AX buf_r_1059__740 (.D(buf_x[1059]), .CK(clock), .Q(buf_r[1059]));
    defparam buf_r_1059__740.GSR = "DISABLED";
    FD1S3AX buf_r_1058__741 (.D(buf_x[1058]), .CK(clock), .Q(buf_r[1058]));
    defparam buf_r_1058__741.GSR = "DISABLED";
    FD1S3AX buf_r_1057__742 (.D(buf_x[1057]), .CK(clock), .Q(buf_r[1057]));
    defparam buf_r_1057__742.GSR = "DISABLED";
    FD1S3AX buf_r_1056__743 (.D(buf_x[1056]), .CK(clock), .Q(buf_r[1056]));
    defparam buf_r_1056__743.GSR = "DISABLED";
    FD1S3AX buf_r_1055__744 (.D(buf_x[1055]), .CK(clock), .Q(buf_r[1055]));
    defparam buf_r_1055__744.GSR = "DISABLED";
    FD1S3AX buf_r_1054__745 (.D(buf_x[1054]), .CK(clock), .Q(buf_r[1054]));
    defparam buf_r_1054__745.GSR = "DISABLED";
    FD1S3AX buf_r_1051__748 (.D(buf_x[1051]), .CK(clock), .Q(buf_r[1051]));
    defparam buf_r_1051__748.GSR = "DISABLED";
    FD1S3AX buf_r_1050__749 (.D(buf_x[1050]), .CK(clock), .Q(buf_r[1050]));
    defparam buf_r_1050__749.GSR = "DISABLED";
    FD1S3AX buf_r_1049__750 (.D(buf_x[1049]), .CK(clock), .Q(buf_r[1049]));
    defparam buf_r_1049__750.GSR = "DISABLED";
    FD1S3AX buf_r_1048__751 (.D(buf_x[1048]), .CK(clock), .Q(buf_r[1048]));
    defparam buf_r_1048__751.GSR = "DISABLED";
    FD1S3AX buf_r_1047__752 (.D(buf_x[1047]), .CK(clock), .Q(buf_r[1047]));
    defparam buf_r_1047__752.GSR = "DISABLED";
    FD1S3AX buf_r_1046__753 (.D(buf_x[1046]), .CK(clock), .Q(buf_r[1046]));
    defparam buf_r_1046__753.GSR = "DISABLED";
    FD1S3AX buf_r_1045__754 (.D(buf_x[1045]), .CK(clock), .Q(buf_r[1045]));
    defparam buf_r_1045__754.GSR = "DISABLED";
    FD1S3AX buf_r_1044__755 (.D(buf_x[1044]), .CK(clock), .Q(buf_r[1044]));
    defparam buf_r_1044__755.GSR = "DISABLED";
    FD1S3AX buf_r_1043__756 (.D(buf_x[1043]), .CK(clock), .Q(buf_r[1043]));
    defparam buf_r_1043__756.GSR = "DISABLED";
    FD1S3AX buf_r_1042__757 (.D(buf_x[1042]), .CK(clock), .Q(buf_r[1042]));
    defparam buf_r_1042__757.GSR = "DISABLED";
    FD1S3AX buf_r_1041__758 (.D(buf_x[1041]), .CK(clock), .Q(buf_r[1041]));
    defparam buf_r_1041__758.GSR = "DISABLED";
    FD1S3AX buf_r_1040__759 (.D(buf_x[1040]), .CK(clock), .Q(buf_r[1040]));
    defparam buf_r_1040__759.GSR = "DISABLED";
    FD1S3AX buf_r_1039__760 (.D(buf_x[1039]), .CK(clock), .Q(buf_r[1039]));
    defparam buf_r_1039__760.GSR = "DISABLED";
    FD1S3AX buf_r_1038__761 (.D(buf_x[1038]), .CK(clock), .Q(buf_r[1038]));
    defparam buf_r_1038__761.GSR = "DISABLED";
    FD1S3AX buf_r_1037__762 (.D(buf_x[1037]), .CK(clock), .Q(buf_r[1037]));
    defparam buf_r_1037__762.GSR = "DISABLED";
    FD1S3AX buf_r_1036__763 (.D(buf_x[1036]), .CK(clock), .Q(buf_r[1036]));
    defparam buf_r_1036__763.GSR = "DISABLED";
    FD1S3AX buf_r_1035__764 (.D(buf_x[1035]), .CK(clock), .Q(buf_r[1035]));
    defparam buf_r_1035__764.GSR = "DISABLED";
    FD1S3AX buf_r_1034__765 (.D(buf_x[1034]), .CK(clock), .Q(buf_r[1034]));
    defparam buf_r_1034__765.GSR = "DISABLED";
    FD1S3AX buf_r_1033__766 (.D(buf_x[1033]), .CK(clock), .Q(buf_r[1033]));
    defparam buf_r_1033__766.GSR = "DISABLED";
    FD1S3AX buf_r_1032__767 (.D(buf_x[1032]), .CK(clock), .Q(buf_r[1032]));
    defparam buf_r_1032__767.GSR = "DISABLED";
    FD1S3AX buf_r_1031__768 (.D(buf_x[1031]), .CK(clock), .Q(buf_r[1031]));
    defparam buf_r_1031__768.GSR = "DISABLED";
    FD1S3AX buf_r_1030__769 (.D(buf_x[1030]), .CK(clock), .Q(buf_r[1030]));
    defparam buf_r_1030__769.GSR = "DISABLED";
    FD1S3AX buf_r_1029__770 (.D(buf_x[1029]), .CK(clock), .Q(buf_r[1029]));
    defparam buf_r_1029__770.GSR = "DISABLED";
    FD1S3AX buf_r_1028__771 (.D(buf_x[1028]), .CK(clock), .Q(buf_r[1028]));
    defparam buf_r_1028__771.GSR = "DISABLED";
    FD1S3AX buf_r_1027__772 (.D(buf_x[1027]), .CK(clock), .Q(buf_r[1027]));
    defparam buf_r_1027__772.GSR = "DISABLED";
    FD1S3AX buf_r_1026__773 (.D(buf_x[1026]), .CK(clock), .Q(buf_r[1026]));
    defparam buf_r_1026__773.GSR = "DISABLED";
    FD1S3AX buf_r_1025__774 (.D(buf_x[1025]), .CK(clock), .Q(buf_r[1025]));
    defparam buf_r_1025__774.GSR = "DISABLED";
    FD1S3AX buf_r_1024__775 (.D(buf_x[1024]), .CK(clock), .Q(buf_r[1024]));
    defparam buf_r_1024__775.GSR = "DISABLED";
    FD1S3AX buf_r_1023__776 (.D(buf_x[1023]), .CK(clock), .Q(buf_x[1490]));
    defparam buf_r_1023__776.GSR = "DISABLED";
    FD1S3AX buf_r_1020__779 (.D(buf_x[1020]), .CK(clock), .Q(buf_r[1020]));
    defparam buf_r_1020__779.GSR = "DISABLED";
    FD1S3AX buf_r_1019__780 (.D(buf_x[1019]), .CK(clock), .Q(buf_r[1019]));
    defparam buf_r_1019__780.GSR = "DISABLED";
    FD1S3AX buf_r_1018__781 (.D(buf_x[1018]), .CK(clock), .Q(buf_r[1018]));
    defparam buf_r_1018__781.GSR = "DISABLED";
    FD1S3AX buf_r_1017__782 (.D(buf_x[1017]), .CK(clock), .Q(buf_r[1017]));
    defparam buf_r_1017__782.GSR = "DISABLED";
    FD1S3AX buf_r_1016__783 (.D(buf_x[1016]), .CK(clock), .Q(buf_r[1016]));
    defparam buf_r_1016__783.GSR = "DISABLED";
    FD1S3AX buf_r_1015__784 (.D(buf_x[1015]), .CK(clock), .Q(buf_r[1015]));
    defparam buf_r_1015__784.GSR = "DISABLED";
    FD1S3AX buf_r_1014__785 (.D(buf_x[1014]), .CK(clock), .Q(buf_r[1014]));
    defparam buf_r_1014__785.GSR = "DISABLED";
    FD1S3AX buf_r_1013__786 (.D(buf_x[1013]), .CK(clock), .Q(buf_r[1013]));
    defparam buf_r_1013__786.GSR = "DISABLED";
    FD1S3AX buf_r_1012__787 (.D(buf_x[1012]), .CK(clock), .Q(buf_r[1012]));
    defparam buf_r_1012__787.GSR = "DISABLED";
    FD1S3AX buf_r_1011__788 (.D(buf_x[1011]), .CK(clock), .Q(buf_r[1011]));
    defparam buf_r_1011__788.GSR = "DISABLED";
    FD1S3AX buf_r_1010__789 (.D(buf_x[1010]), .CK(clock), .Q(buf_r[1010]));
    defparam buf_r_1010__789.GSR = "DISABLED";
    FD1S3AX buf_r_1009__790 (.D(buf_x[1009]), .CK(clock), .Q(buf_r[1009]));
    defparam buf_r_1009__790.GSR = "DISABLED";
    FD1S3AX buf_r_1008__791 (.D(buf_x[1008]), .CK(clock), .Q(buf_r[1008]));
    defparam buf_r_1008__791.GSR = "DISABLED";
    FD1S3AX buf_r_1007__792 (.D(buf_x[1007]), .CK(clock), .Q(buf_r[1007]));
    defparam buf_r_1007__792.GSR = "DISABLED";
    FD1S3AX buf_r_1006__793 (.D(buf_x[1006]), .CK(clock), .Q(buf_r[1006]));
    defparam buf_r_1006__793.GSR = "DISABLED";
    FD1S3AX buf_r_1005__794 (.D(buf_x[1005]), .CK(clock), .Q(buf_r[1005]));
    defparam buf_r_1005__794.GSR = "DISABLED";
    FD1S3AX buf_r_1004__795 (.D(buf_x[1004]), .CK(clock), .Q(buf_r[1004]));
    defparam buf_r_1004__795.GSR = "DISABLED";
    FD1S3AX buf_r_1003__796 (.D(buf_x[1003]), .CK(clock), .Q(buf_r[1003]));
    defparam buf_r_1003__796.GSR = "DISABLED";
    FD1S3AX buf_r_1002__797 (.D(buf_x[1002]), .CK(clock), .Q(buf_r[1002]));
    defparam buf_r_1002__797.GSR = "DISABLED";
    FD1S3AX buf_r_1001__798 (.D(buf_x[1001]), .CK(clock), .Q(buf_r[1001]));
    defparam buf_r_1001__798.GSR = "DISABLED";
    FD1S3AX buf_r_1000__799 (.D(buf_x[1000]), .CK(clock), .Q(buf_r[1000]));
    defparam buf_r_1000__799.GSR = "DISABLED";
    FD1S3AX buf_r_999__800 (.D(buf_x[999]), .CK(clock), .Q(buf_r[999]));
    defparam buf_r_999__800.GSR = "DISABLED";
    FD1S3AX buf_r_998__801 (.D(buf_x[998]), .CK(clock), .Q(buf_r[998]));
    defparam buf_r_998__801.GSR = "DISABLED";
    FD1S3AX buf_r_997__802 (.D(buf_x[997]), .CK(clock), .Q(buf_r[997]));
    defparam buf_r_997__802.GSR = "DISABLED";
    FD1S3AX buf_r_996__803 (.D(buf_x[996]), .CK(clock), .Q(buf_r[996]));
    defparam buf_r_996__803.GSR = "DISABLED";
    FD1S3AX buf_r_995__804 (.D(buf_x[995]), .CK(clock), .Q(buf_r[995]));
    defparam buf_r_995__804.GSR = "DISABLED";
    FD1S3AX buf_r_994__805 (.D(buf_x[994]), .CK(clock), .Q(buf_r[994]));
    defparam buf_r_994__805.GSR = "DISABLED";
    FD1S3AX buf_r_993__806 (.D(buf_x[993]), .CK(clock), .Q(buf_r[993]));
    defparam buf_r_993__806.GSR = "DISABLED";
    FD1S3AX buf_r_992__807 (.D(buf_x[992]), .CK(clock), .Q(buf_r[992]));
    defparam buf_r_992__807.GSR = "DISABLED";
    FD1S3AX buf_r_989__810 (.D(buf_x[989]), .CK(clock), .Q(buf_r[989]));
    defparam buf_r_989__810.GSR = "DISABLED";
    FD1S3AX buf_r_988__811 (.D(buf_x[988]), .CK(clock), .Q(buf_r[988]));
    defparam buf_r_988__811.GSR = "DISABLED";
    FD1S3AX buf_r_987__812 (.D(buf_x[987]), .CK(clock), .Q(buf_r[987]));
    defparam buf_r_987__812.GSR = "DISABLED";
    FD1S3AX buf_r_986__813 (.D(buf_x[986]), .CK(clock), .Q(buf_r[986]));
    defparam buf_r_986__813.GSR = "DISABLED";
    FD1S3AX buf_r_985__814 (.D(buf_x[985]), .CK(clock), .Q(buf_r[985]));
    defparam buf_r_985__814.GSR = "DISABLED";
    FD1S3AX buf_r_984__815 (.D(buf_x[984]), .CK(clock), .Q(buf_r[984]));
    defparam buf_r_984__815.GSR = "DISABLED";
    FD1S3AX buf_r_983__816 (.D(buf_x[983]), .CK(clock), .Q(buf_r[983]));
    defparam buf_r_983__816.GSR = "DISABLED";
    FD1S3AX buf_r_982__817 (.D(buf_x[982]), .CK(clock), .Q(buf_r[982]));
    defparam buf_r_982__817.GSR = "DISABLED";
    FD1S3AX buf_r_981__818 (.D(buf_x[981]), .CK(clock), .Q(buf_r[981]));
    defparam buf_r_981__818.GSR = "DISABLED";
    FD1S3AX buf_r_980__819 (.D(buf_x[980]), .CK(clock), .Q(buf_r[980]));
    defparam buf_r_980__819.GSR = "DISABLED";
    FD1S3AX buf_r_979__820 (.D(buf_x[979]), .CK(clock), .Q(buf_r[979]));
    defparam buf_r_979__820.GSR = "DISABLED";
    FD1S3AX buf_r_978__821 (.D(buf_x[978]), .CK(clock), .Q(buf_r[978]));
    defparam buf_r_978__821.GSR = "DISABLED";
    FD1S3AX buf_r_977__822 (.D(buf_x[977]), .CK(clock), .Q(buf_r[977]));
    defparam buf_r_977__822.GSR = "DISABLED";
    FD1S3AX buf_r_976__823 (.D(buf_x[976]), .CK(clock), .Q(buf_r[976]));
    defparam buf_r_976__823.GSR = "DISABLED";
    FD1S3AX buf_r_975__824 (.D(buf_x[975]), .CK(clock), .Q(buf_r[975]));
    defparam buf_r_975__824.GSR = "DISABLED";
    FD1S3AX buf_r_974__825 (.D(buf_x[974]), .CK(clock), .Q(buf_r[974]));
    defparam buf_r_974__825.GSR = "DISABLED";
    FD1S3AX buf_r_973__826 (.D(buf_x[973]), .CK(clock), .Q(buf_r[973]));
    defparam buf_r_973__826.GSR = "DISABLED";
    FD1S3AX buf_r_972__827 (.D(buf_x[972]), .CK(clock), .Q(buf_r[972]));
    defparam buf_r_972__827.GSR = "DISABLED";
    FD1S3AX buf_r_971__828 (.D(buf_x[971]), .CK(clock), .Q(buf_r[971]));
    defparam buf_r_971__828.GSR = "DISABLED";
    FD1S3AX buf_r_970__829 (.D(buf_x[970]), .CK(clock), .Q(buf_r[970]));
    defparam buf_r_970__829.GSR = "DISABLED";
    FD1S3AX buf_r_969__830 (.D(buf_x[969]), .CK(clock), .Q(buf_r[969]));
    defparam buf_r_969__830.GSR = "DISABLED";
    FD1S3AX buf_r_968__831 (.D(buf_x[968]), .CK(clock), .Q(buf_r[968]));
    defparam buf_r_968__831.GSR = "DISABLED";
    FD1S3AX buf_r_967__832 (.D(buf_x[967]), .CK(clock), .Q(buf_r[967]));
    defparam buf_r_967__832.GSR = "DISABLED";
    FD1S3AX buf_r_966__833 (.D(buf_x[966]), .CK(clock), .Q(buf_r[966]));
    defparam buf_r_966__833.GSR = "DISABLED";
    FD1S3AX buf_r_965__834 (.D(buf_x[965]), .CK(clock), .Q(buf_r[965]));
    defparam buf_r_965__834.GSR = "DISABLED";
    FD1S3AX buf_r_964__835 (.D(buf_x[964]), .CK(clock), .Q(buf_r[964]));
    defparam buf_r_964__835.GSR = "DISABLED";
    FD1S3AX buf_r_963__836 (.D(buf_x[963]), .CK(clock), .Q(buf_r[963]));
    defparam buf_r_963__836.GSR = "DISABLED";
    FD1S3AX buf_r_962__837 (.D(buf_x[962]), .CK(clock), .Q(buf_r[962]));
    defparam buf_r_962__837.GSR = "DISABLED";
    FD1S3AX buf_r_1827__843 (.D(buf_x[1827]), .CK(clock), .Q(buf_x[1946]));
    defparam buf_r_1827__843.GSR = "DISABLED";
    FD1S3AX buf_r_1826__844 (.D(buf_x[1826]), .CK(clock), .Q(buf_x[1945]));
    defparam buf_r_1826__844.GSR = "DISABLED";
    FD1S3AX buf_r_1825__845 (.D(buf_x[1825]), .CK(clock), .Q(buf_x[1944]));
    defparam buf_r_1825__845.GSR = "DISABLED";
    FD1S3AX buf_r_1824__846 (.D(buf_x[1824]), .CK(clock), .Q(buf_x[1943]));
    defparam buf_r_1824__846.GSR = "DISABLED";
    FD1S3AX buf_r_1823__847 (.D(buf_x[1823]), .CK(clock), .Q(buf_x[1942]));
    defparam buf_r_1823__847.GSR = "DISABLED";
    FD1S3AX buf_r_1822__848 (.D(buf_x[1822]), .CK(clock), .Q(buf_x[1941]));
    defparam buf_r_1822__848.GSR = "DISABLED";
    FD1S3AX buf_r_1821__849 (.D(buf_x[1821]), .CK(clock), .Q(buf_x[1940]));
    defparam buf_r_1821__849.GSR = "DISABLED";
    FD1S3AX buf_r_1820__850 (.D(buf_x[1820]), .CK(clock), .Q(buf_x[1939]));
    defparam buf_r_1820__850.GSR = "DISABLED";
    FD1S3AX buf_r_1819__851 (.D(buf_x[1819]), .CK(clock), .Q(buf_x[1938]));
    defparam buf_r_1819__851.GSR = "DISABLED";
    FD1S3AX buf_r_1818__852 (.D(buf_x[1818]), .CK(clock), .Q(buf_x[1937]));
    defparam buf_r_1818__852.GSR = "DISABLED";
    FD1S3AX buf_r_1817__853 (.D(buf_x[1817]), .CK(clock), .Q(buf_x[1936]));
    defparam buf_r_1817__853.GSR = "DISABLED";
    FD1S3AX buf_r_1816__854 (.D(buf_x[1816]), .CK(clock), .Q(buf_x[1935]));
    defparam buf_r_1816__854.GSR = "DISABLED";
    FD1S3AX buf_r_1815__855 (.D(buf_x[1815]), .CK(clock), .Q(buf_x[1934]));
    defparam buf_r_1815__855.GSR = "DISABLED";
    FD1S3AX buf_r_1814__856 (.D(buf_x[1814]), .CK(clock), .Q(buf_x[1933]));
    defparam buf_r_1814__856.GSR = "DISABLED";
    FD1S3AX buf_r_1813__857 (.D(buf_x[1813]), .CK(clock), .Q(buf_x[1932]));
    defparam buf_r_1813__857.GSR = "DISABLED";
    FD1S3AX buf_r_1812__858 (.D(buf_x[1812]), .CK(clock), .Q(buf_x[1931]));
    defparam buf_r_1812__858.GSR = "DISABLED";
    FD1S3AX buf_r_1811__859 (.D(buf_x[1811]), .CK(clock), .Q(buf_x[1930]));
    defparam buf_r_1811__859.GSR = "DISABLED";
    FD1S3AX buf_r_1810__860 (.D(buf_x[1810]), .CK(clock), .Q(buf_x[1929]));
    defparam buf_r_1810__860.GSR = "DISABLED";
    FD1S3AX buf_r_1809__861 (.D(buf_x[1809]), .CK(clock), .Q(buf_x[1928]));
    defparam buf_r_1809__861.GSR = "DISABLED";
    FD1S3AX buf_r_1808__862 (.D(buf_x[1808]), .CK(clock), .Q(buf_x[1927]));
    defparam buf_r_1808__862.GSR = "DISABLED";
    FD1S3AX buf_r_1807__863 (.D(buf_x[1807]), .CK(clock), .Q(buf_x[1926]));
    defparam buf_r_1807__863.GSR = "DISABLED";
    FD1S3AX buf_r_1806__864 (.D(buf_x[1806]), .CK(clock), .Q(buf_x[1925]));
    defparam buf_r_1806__864.GSR = "DISABLED";
    FD1S3AX buf_r_1805__865 (.D(buf_x[1805]), .CK(clock), .Q(buf_x[1924]));
    defparam buf_r_1805__865.GSR = "DISABLED";
    FD1S3AX buf_r_1804__866 (.D(buf_x[1804]), .CK(clock), .Q(buf_x[1923]));
    defparam buf_r_1804__866.GSR = "DISABLED";
    FD1S3AX buf_r_1803__867 (.D(buf_x[1803]), .CK(clock), .Q(buf_x[1922]));
    defparam buf_r_1803__867.GSR = "DISABLED";
    FD1S3AX buf_r_1802__868 (.D(buf_x[1802]), .CK(clock), .Q(buf_x[1921]));
    defparam buf_r_1802__868.GSR = "DISABLED";
    FD1S3AX buf_r_1801__869 (.D(buf_x[1801]), .CK(clock), .Q(buf_x[1920]));
    defparam buf_r_1801__869.GSR = "DISABLED";
    FD1S3AX buf_r_1800__870 (.D(buf_x[1800]), .CK(clock), .Q(buf_x[1919]));
    defparam buf_r_1800__870.GSR = "DISABLED";
    FD1S3AX buf_r_1799__871 (.D(buf_x[1799]), .CK(clock), .Q(buf_x[1918]));
    defparam buf_r_1799__871.GSR = "DISABLED";
    FD1S3AX buf_r_1798__872 (.D(buf_x[1798]), .CK(clock), .Q(buf_x[1917]));
    defparam buf_r_1798__872.GSR = "DISABLED";
    FD1S3AX buf_r_1797__873 (.D(buf_x[1797]), .CK(clock), .Q(buf_x[1916]));
    defparam buf_r_1797__873.GSR = "DISABLED";
    FD1S3AX buf_r_1796__874 (.D(buf_x[1796]), .CK(clock), .Q(buf_x[1915]));
    defparam buf_r_1796__874.GSR = "DISABLED";
    FD1S3AX buf_r_1795__875 (.D(buf_x[1795]), .CK(clock), .Q(buf_x[1914]));
    defparam buf_r_1795__875.GSR = "DISABLED";
    FD1S3AX buf_r_1794__876 (.D(buf_x[1794]), .CK(clock), .Q(buf_x[1913]));
    defparam buf_r_1794__876.GSR = "DISABLED";
    FD1S3AX buf_r_1793__877 (.D(buf_x[1793]), .CK(clock), .Q(buf_r[1793]));
    defparam buf_r_1793__877.GSR = "DISABLED";
    FD1S3AX buf_r_1792__878 (.D(buf_x[1792]), .CK(clock), .Q(buf_r[1792]));
    defparam buf_r_1792__878.GSR = "DISABLED";
    FD1S3AX buf_r_1791__879 (.D(buf_x[1791]), .CK(clock), .Q(buf_r[1791]));
    defparam buf_r_1791__879.GSR = "DISABLED";
    FD1S3AX buf_r_1790__880 (.D(buf_x[1790]), .CK(clock), .Q(buf_r[1790]));
    defparam buf_r_1790__880.GSR = "DISABLED";
    FD1S3AX buf_r_1789__881 (.D(buf_x[1789]), .CK(clock), .Q(buf_r[1789]));
    defparam buf_r_1789__881.GSR = "DISABLED";
    FD1S3AX buf_r_1788__882 (.D(buf_x[1788]), .CK(clock), .Q(buf_r[1788]));
    defparam buf_r_1788__882.GSR = "DISABLED";
    FD1S3AX buf_r_1787__883 (.D(buf_x[1787]), .CK(clock), .Q(buf_r[1787]));
    defparam buf_r_1787__883.GSR = "DISABLED";
    FD1S3AX buf_r_1786__884 (.D(buf_x[1786]), .CK(clock), .Q(buf_r[1786]));
    defparam buf_r_1786__884.GSR = "DISABLED";
    FD1S3AX buf_r_1785__885 (.D(buf_x[1785]), .CK(clock), .Q(buf_r[1785]));
    defparam buf_r_1785__885.GSR = "DISABLED";
    FD1S3AX buf_r_1784__886 (.D(buf_x[1784]), .CK(clock), .Q(buf_r[1784]));
    defparam buf_r_1784__886.GSR = "DISABLED";
    FD1S3AX buf_r_1783__887 (.D(buf_x[1783]), .CK(clock), .Q(buf_r[1783]));
    defparam buf_r_1783__887.GSR = "DISABLED";
    FD1S3AX buf_r_1782__888 (.D(buf_x[1782]), .CK(clock), .Q(buf_r[1782]));
    defparam buf_r_1782__888.GSR = "DISABLED";
    FD1S3AX buf_r_1781__889 (.D(buf_x[1781]), .CK(clock), .Q(buf_r[1781]));
    defparam buf_r_1781__889.GSR = "DISABLED";
    FD1S3AX buf_r_1780__890 (.D(buf_x[1780]), .CK(clock), .Q(buf_r[1780]));
    defparam buf_r_1780__890.GSR = "DISABLED";
    FD1S3AX buf_r_1779__891 (.D(buf_x[1779]), .CK(clock), .Q(buf_r[1779]));
    defparam buf_r_1779__891.GSR = "DISABLED";
    FD1S3AX buf_r_1778__892 (.D(buf_x[1778]), .CK(clock), .Q(buf_r[1778]));
    defparam buf_r_1778__892.GSR = "DISABLED";
    FD1S3AX buf_r_1777__893 (.D(buf_x[1777]), .CK(clock), .Q(buf_r[1777]));
    defparam buf_r_1777__893.GSR = "DISABLED";
    FD1S3AX buf_r_1776__894 (.D(buf_x[1776]), .CK(clock), .Q(buf_r[1776]));
    defparam buf_r_1776__894.GSR = "DISABLED";
    FD1S3AX buf_r_1775__895 (.D(buf_x[1775]), .CK(clock), .Q(buf_r[1775]));
    defparam buf_r_1775__895.GSR = "DISABLED";
    FD1S3AX buf_r_1774__896 (.D(buf_x[1774]), .CK(clock), .Q(buf_r[1774]));
    defparam buf_r_1774__896.GSR = "DISABLED";
    FD1S3AX buf_r_1773__897 (.D(buf_x[1773]), .CK(clock), .Q(buf_r[1773]));
    defparam buf_r_1773__897.GSR = "DISABLED";
    FD1S3AX buf_r_1772__898 (.D(buf_x[1772]), .CK(clock), .Q(buf_r[1772]));
    defparam buf_r_1772__898.GSR = "DISABLED";
    FD1S3AX buf_r_1771__899 (.D(buf_x[1771]), .CK(clock), .Q(buf_r[1771]));
    defparam buf_r_1771__899.GSR = "DISABLED";
    FD1S3AX buf_r_1770__900 (.D(buf_x[1770]), .CK(clock), .Q(buf_r[1770]));
    defparam buf_r_1770__900.GSR = "DISABLED";
    FD1S3AX buf_r_1769__901 (.D(buf_x[1769]), .CK(clock), .Q(buf_r[1769]));
    defparam buf_r_1769__901.GSR = "DISABLED";
    FD1S3AX buf_r_1768__902 (.D(buf_x[1768]), .CK(clock), .Q(buf_r[1768]));
    defparam buf_r_1768__902.GSR = "DISABLED";
    FD1S3AX buf_r_1767__903 (.D(buf_x[1767]), .CK(clock), .Q(buf_r[1767]));
    defparam buf_r_1767__903.GSR = "DISABLED";
    FD1S3AX buf_r_1766__904 (.D(buf_x[1766]), .CK(clock), .Q(buf_r[1766]));
    defparam buf_r_1766__904.GSR = "DISABLED";
    FD1S3AX buf_r_1765__905 (.D(buf_x[1765]), .CK(clock), .Q(buf_r[1765]));
    defparam buf_r_1765__905.GSR = "DISABLED";
    FD1S3AX buf_r_1764__906 (.D(buf_x[1764]), .CK(clock), .Q(buf_r[1764]));
    defparam buf_r_1764__906.GSR = "DISABLED";
    FD1S3AX buf_r_1763__907 (.D(buf_x[1763]), .CK(clock), .Q(buf_r[1763]));
    defparam buf_r_1763__907.GSR = "DISABLED";
    FD1S3AX buf_r_1762__908 (.D(buf_x[1762]), .CK(clock), .Q(buf_r[1762]));
    defparam buf_r_1762__908.GSR = "DISABLED";
    FD1S3AX buf_r_1761__909 (.D(buf_x[1761]), .CK(clock), .Q(buf_r[1761]));
    defparam buf_r_1761__909.GSR = "DISABLED";
    FD1S3AX buf_r_1760__910 (.D(buf_x[1760]), .CK(clock), .Q(buf_r[1760]));
    defparam buf_r_1760__910.GSR = "DISABLED";
    FD1S3AX buf_r_1759__911 (.D(buf_x[1759]), .CK(clock), .Q(buf_r[1759]));
    defparam buf_r_1759__911.GSR = "DISABLED";
    FD1S3AX buf_r_1758__912 (.D(buf_x[1758]), .CK(clock), .Q(buf_r[1758]));
    defparam buf_r_1758__912.GSR = "DISABLED";
    FD1S3AX buf_r_1757__913 (.D(buf_x[1757]), .CK(clock), .Q(buf_r[1757]));
    defparam buf_r_1757__913.GSR = "DISABLED";
    FD1S3AX buf_r_1756__914 (.D(buf_x[1756]), .CK(clock), .Q(buf_r[1756]));
    defparam buf_r_1756__914.GSR = "DISABLED";
    FD1S3AX buf_r_1755__915 (.D(buf_x[1755]), .CK(clock), .Q(buf_r[1755]));
    defparam buf_r_1755__915.GSR = "DISABLED";
    FD1S3AX buf_r_1754__916 (.D(buf_x[1754]), .CK(clock), .Q(buf_r[1754]));
    defparam buf_r_1754__916.GSR = "DISABLED";
    FD1S3AX buf_r_1753__917 (.D(buf_x[1753]), .CK(clock), .Q(buf_r[1753]));
    defparam buf_r_1753__917.GSR = "DISABLED";
    FD1S3AX buf_r_1752__918 (.D(buf_x[1752]), .CK(clock), .Q(buf_r[1752]));
    defparam buf_r_1752__918.GSR = "DISABLED";
    FD1S3AX buf_r_1751__919 (.D(buf_x[1751]), .CK(clock), .Q(buf_r[1751]));
    defparam buf_r_1751__919.GSR = "DISABLED";
    FD1S3AX buf_r_1750__920 (.D(buf_x[1750]), .CK(clock), .Q(buf_r[1750]));
    defparam buf_r_1750__920.GSR = "DISABLED";
    FD1S3AX buf_r_1749__921 (.D(buf_x[1749]), .CK(clock), .Q(buf_r[1749]));
    defparam buf_r_1749__921.GSR = "DISABLED";
    FD1S3AX buf_r_1748__922 (.D(buf_x[1748]), .CK(clock), .Q(buf_r[1748]));
    defparam buf_r_1748__922.GSR = "DISABLED";
    FD1S3AX buf_r_1747__923 (.D(buf_x[1747]), .CK(clock), .Q(buf_r[1747]));
    defparam buf_r_1747__923.GSR = "DISABLED";
    FD1S3AX buf_r_1746__924 (.D(buf_x[1746]), .CK(clock), .Q(buf_r[1746]));
    defparam buf_r_1746__924.GSR = "DISABLED";
    FD1S3AX buf_r_1745__925 (.D(buf_x[1745]), .CK(clock), .Q(buf_r[1745]));
    defparam buf_r_1745__925.GSR = "DISABLED";
    FD1S3AX buf_r_1744__926 (.D(buf_x[1744]), .CK(clock), .Q(buf_r[1744]));
    defparam buf_r_1744__926.GSR = "DISABLED";
    FD1S3AX buf_r_1743__927 (.D(buf_x[1743]), .CK(clock), .Q(buf_r[1743]));
    defparam buf_r_1743__927.GSR = "DISABLED";
    FD1S3AX buf_r_1742__928 (.D(buf_x[1742]), .CK(clock), .Q(buf_r[1742]));
    defparam buf_r_1742__928.GSR = "DISABLED";
    FD1S3AX buf_r_1741__929 (.D(buf_x[1741]), .CK(clock), .Q(buf_r[1741]));
    defparam buf_r_1741__929.GSR = "DISABLED";
    FD1S3AX buf_r_1740__930 (.D(buf_x[1740]), .CK(clock), .Q(buf_r[1740]));
    defparam buf_r_1740__930.GSR = "DISABLED";
    FD1S3AX buf_r_1739__931 (.D(buf_x[1739]), .CK(clock), .Q(buf_r[1739]));
    defparam buf_r_1739__931.GSR = "DISABLED";
    FD1S3AX buf_r_1738__932 (.D(buf_x[1738]), .CK(clock), .Q(buf_r[1738]));
    defparam buf_r_1738__932.GSR = "DISABLED";
    FD1S3AX buf_r_1737__933 (.D(buf_x[1737]), .CK(clock), .Q(buf_r[1737]));
    defparam buf_r_1737__933.GSR = "DISABLED";
    FD1S3AX buf_r_1736__934 (.D(buf_x[1736]), .CK(clock), .Q(buf_r[1736]));
    defparam buf_r_1736__934.GSR = "DISABLED";
    FD1S3AX buf_r_1735__935 (.D(buf_x[1735]), .CK(clock), .Q(buf_r[1735]));
    defparam buf_r_1735__935.GSR = "DISABLED";
    FD1S3AX buf_r_1734__936 (.D(buf_x[1734]), .CK(clock), .Q(buf_r[1734]));
    defparam buf_r_1734__936.GSR = "DISABLED";
    FD1S3AX buf_r_1733__937 (.D(buf_x[1733]), .CK(clock), .Q(buf_r[1733]));
    defparam buf_r_1733__937.GSR = "DISABLED";
    FD1S3AX buf_r_1732__938 (.D(buf_x[1732]), .CK(clock), .Q(buf_r[1732]));
    defparam buf_r_1732__938.GSR = "DISABLED";
    FD1S3AX buf_r_1731__939 (.D(buf_x[1731]), .CK(clock), .Q(buf_r[1731]));
    defparam buf_r_1731__939.GSR = "DISABLED";
    FD1S3AX buf_r_1730__940 (.D(buf_x[1730]), .CK(clock), .Q(buf_r[1730]));
    defparam buf_r_1730__940.GSR = "DISABLED";
    FD1S3AX buf_r_1729__941 (.D(buf_x[1729]), .CK(clock), .Q(buf_r[1729]));
    defparam buf_r_1729__941.GSR = "DISABLED";
    FD1S3AX buf_r_1728__942 (.D(buf_x[1728]), .CK(clock), .Q(buf_r[1728]));
    defparam buf_r_1728__942.GSR = "DISABLED";
    CCU2D add_4611_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[16]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[15]), .B1(nZ0_d2[16]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[17]), .CIN(n61965), .COUT(n61966), .S0(buf_x[1222]), 
          .S1(buf_x[1223]));
    defparam add_4611_15.INIT0 = 16'h7888;
    defparam add_4611_15.INIT1 = 16'h7888;
    defparam add_4611_15.INJECT1_0 = "NO";
    defparam add_4611_15.INJECT1_1 = "NO";
    CCU2D add_4611_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[16]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[13]), .B1(nZ0_d2[16]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[17]), .CIN(n61964), .COUT(n61965), .S0(buf_x[1220]), 
          .S1(buf_x[1221]));
    defparam add_4611_13.INIT0 = 16'h7888;
    defparam add_4611_13.INIT1 = 16'h7888;
    defparam add_4611_13.INJECT1_0 = "NO";
    defparam add_4611_13.INJECT1_1 = "NO";
    CCU2D add_4611_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[16]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[11]), .B1(nZ0_d2[16]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[17]), .CIN(n61963), .COUT(n61964), .S0(buf_x[1218]), 
          .S1(buf_x[1219]));
    defparam add_4611_11.INIT0 = 16'h7888;
    defparam add_4611_11.INIT1 = 16'h7888;
    defparam add_4611_11.INJECT1_0 = "NO";
    defparam add_4611_11.INJECT1_1 = "NO";
    CCU2D add_4611_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[16]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[9]), .B1(nZ0_d2[16]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[17]), .CIN(n61962), .COUT(n61963), .S0(buf_x[1216]), 
          .S1(buf_x[1217]));
    defparam add_4611_9.INIT0 = 16'h7888;
    defparam add_4611_9.INIT1 = 16'h7888;
    defparam add_4611_9.INJECT1_0 = "NO";
    defparam add_4611_9.INJECT1_1 = "NO";
    CCU2D add_4611_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[16]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[7]), .B1(nZ0_d2[16]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[17]), .CIN(n61961), .COUT(n61962), .S0(buf_x[1214]), 
          .S1(buf_x[1215]));
    defparam add_4611_7.INIT0 = 16'h7888;
    defparam add_4611_7.INIT1 = 16'h7888;
    defparam add_4611_7.INJECT1_0 = "NO";
    defparam add_4611_7.INJECT1_1 = "NO";
    CCU2D add_4611_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[16]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[5]), .B1(nZ0_d2[16]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[17]), .CIN(n61960), .COUT(n61961), .S0(buf_x[1212]), 
          .S1(buf_x[1213]));
    defparam add_4611_5.INIT0 = 16'h7888;
    defparam add_4611_5.INIT1 = 16'h7888;
    defparam add_4611_5.INJECT1_0 = "NO";
    defparam add_4611_5.INJECT1_1 = "NO";
    CCU2D add_4611_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[16]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[17]), .A1(nEY1_d2[3]), .B1(nZ0_d2[16]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[17]), .CIN(n61959), .COUT(n61960), .S0(buf_x[1210]), 
          .S1(buf_x[1211]));
    defparam add_4611_3.INIT0 = 16'h7888;
    defparam add_4611_3.INIT1 = 16'h7888;
    defparam add_4611_3.INJECT1_0 = "NO";
    defparam add_4611_3.INJECT1_1 = "NO";
    CCU2D add_4611_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[16]), .C1(nEY1_d2[0]), .D1(nZ0_d2[17]), 
          .COUT(n61959), .S1(buf_x[1209]));
    defparam add_4611_1.INIT0 = 16'hF000;
    defparam add_4611_1.INIT1 = 16'h7888;
    defparam add_4611_1.INJECT1_0 = "NO";
    defparam add_4611_1.INJECT1_1 = "NO";
    CCU2D add_4610_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[15]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61958), .S0(buf_x[1205]), .S1(buf_x[1206]));
    defparam add_4610_29.INIT0 = 16'h7888;
    defparam add_4610_29.INIT1 = 16'h0000;
    defparam add_4610_29.INJECT1_0 = "NO";
    defparam add_4610_29.INJECT1_1 = "NO";
    CCU2D add_4610_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[14]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[27]), .B1(nZ0_d2[14]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[15]), .CIN(n61957), .COUT(n61958), .S0(buf_x[1203]), 
          .S1(buf_x[1204]));
    defparam add_4610_27.INIT0 = 16'h7888;
    defparam add_4610_27.INIT1 = 16'h7888;
    defparam add_4610_27.INJECT1_0 = "NO";
    defparam add_4610_27.INJECT1_1 = "NO";
    CCU2D add_4610_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[14]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[25]), .B1(nZ0_d2[14]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[15]), .CIN(n61956), .COUT(n61957), .S0(buf_x[1201]), 
          .S1(buf_x[1202]));
    defparam add_4610_25.INIT0 = 16'h7888;
    defparam add_4610_25.INIT1 = 16'h7888;
    defparam add_4610_25.INJECT1_0 = "NO";
    defparam add_4610_25.INJECT1_1 = "NO";
    CCU2D add_4610_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[14]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[23]), .B1(nZ0_d2[14]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[15]), .CIN(n61955), .COUT(n61956), .S0(buf_x[1199]), 
          .S1(buf_x[1200]));
    defparam add_4610_23.INIT0 = 16'h7888;
    defparam add_4610_23.INIT1 = 16'h7888;
    defparam add_4610_23.INJECT1_0 = "NO";
    defparam add_4610_23.INJECT1_1 = "NO";
    CCU2D add_4610_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[14]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[21]), .B1(nZ0_d2[14]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[15]), .CIN(n61954), .COUT(n61955), .S0(buf_x[1197]), 
          .S1(buf_x[1198]));
    defparam add_4610_21.INIT0 = 16'h7888;
    defparam add_4610_21.INIT1 = 16'h7888;
    defparam add_4610_21.INJECT1_0 = "NO";
    defparam add_4610_21.INJECT1_1 = "NO";
    CCU2D add_4610_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[14]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[19]), .B1(nZ0_d2[14]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[15]), .CIN(n61953), .COUT(n61954), .S0(buf_x[1195]), 
          .S1(buf_x[1196]));
    defparam add_4610_19.INIT0 = 16'h7888;
    defparam add_4610_19.INIT1 = 16'h7888;
    defparam add_4610_19.INJECT1_0 = "NO";
    defparam add_4610_19.INJECT1_1 = "NO";
    CCU2D add_4610_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[14]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[17]), .B1(nZ0_d2[14]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[15]), .CIN(n61952), .COUT(n61953), .S0(buf_x[1193]), 
          .S1(buf_x[1194]));
    defparam add_4610_17.INIT0 = 16'h7888;
    defparam add_4610_17.INIT1 = 16'h7888;
    defparam add_4610_17.INJECT1_0 = "NO";
    defparam add_4610_17.INJECT1_1 = "NO";
    CCU2D add_4610_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[14]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[15]), .B1(nZ0_d2[14]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[15]), .CIN(n61951), .COUT(n61952), .S0(buf_x[1191]), 
          .S1(buf_x[1192]));
    defparam add_4610_15.INIT0 = 16'h7888;
    defparam add_4610_15.INIT1 = 16'h7888;
    defparam add_4610_15.INJECT1_0 = "NO";
    defparam add_4610_15.INJECT1_1 = "NO";
    CCU2D add_4610_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[14]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[13]), .B1(nZ0_d2[14]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[15]), .CIN(n61950), .COUT(n61951), .S0(buf_x[1189]), 
          .S1(buf_x[1190]));
    defparam add_4610_13.INIT0 = 16'h7888;
    defparam add_4610_13.INIT1 = 16'h7888;
    defparam add_4610_13.INJECT1_0 = "NO";
    defparam add_4610_13.INJECT1_1 = "NO";
    CCU2D add_4610_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[14]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[11]), .B1(nZ0_d2[14]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[15]), .CIN(n61949), .COUT(n61950), .S0(buf_x[1187]), 
          .S1(buf_x[1188]));
    defparam add_4610_11.INIT0 = 16'h7888;
    defparam add_4610_11.INIT1 = 16'h7888;
    defparam add_4610_11.INJECT1_0 = "NO";
    defparam add_4610_11.INJECT1_1 = "NO";
    CCU2D add_4610_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[14]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[9]), .B1(nZ0_d2[14]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[15]), .CIN(n61948), .COUT(n61949), .S0(buf_x[1185]), 
          .S1(buf_x[1186]));
    defparam add_4610_9.INIT0 = 16'h7888;
    defparam add_4610_9.INIT1 = 16'h7888;
    defparam add_4610_9.INJECT1_0 = "NO";
    defparam add_4610_9.INJECT1_1 = "NO";
    CCU2D add_4610_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[14]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[7]), .B1(nZ0_d2[14]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[15]), .CIN(n61947), .COUT(n61948), .S0(buf_x[1183]), 
          .S1(buf_x[1184]));
    defparam add_4610_7.INIT0 = 16'h7888;
    defparam add_4610_7.INIT1 = 16'h7888;
    defparam add_4610_7.INJECT1_0 = "NO";
    defparam add_4610_7.INJECT1_1 = "NO";
    CCU2D add_4610_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[14]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[5]), .B1(nZ0_d2[14]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[15]), .CIN(n61946), .COUT(n61947), .S0(buf_x[1181]), 
          .S1(buf_x[1182]));
    defparam add_4610_5.INIT0 = 16'h7888;
    defparam add_4610_5.INIT1 = 16'h7888;
    defparam add_4610_5.INJECT1_0 = "NO";
    defparam add_4610_5.INJECT1_1 = "NO";
    CCU2D add_4610_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[14]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[15]), .A1(nEY1_d2[3]), .B1(nZ0_d2[14]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[15]), .CIN(n61945), .COUT(n61946), .S0(buf_x[1179]), 
          .S1(buf_x[1180]));
    defparam add_4610_3.INIT0 = 16'h7888;
    defparam add_4610_3.INIT1 = 16'h7888;
    defparam add_4610_3.INJECT1_0 = "NO";
    defparam add_4610_3.INJECT1_1 = "NO";
    CCU2D add_4610_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[14]), .C1(nEY1_d2[0]), .D1(nZ0_d2[15]), 
          .COUT(n61945), .S1(buf_x[1178]));
    defparam add_4610_1.INIT0 = 16'hF000;
    defparam add_4610_1.INIT1 = 16'h7888;
    defparam add_4610_1.INJECT1_0 = "NO";
    defparam add_4610_1.INJECT1_1 = "NO";
    CCU2D add_4609_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[13]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61944), .S0(buf_x[1174]), .S1(buf_x[1175]));
    defparam add_4609_29.INIT0 = 16'h7888;
    defparam add_4609_29.INIT1 = 16'h0000;
    defparam add_4609_29.INJECT1_0 = "NO";
    defparam add_4609_29.INJECT1_1 = "NO";
    CCU2D add_4609_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[12]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[27]), .B1(nZ0_d2[12]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[13]), .CIN(n61943), .COUT(n61944), .S0(buf_x[1172]), 
          .S1(buf_x[1173]));
    defparam add_4609_27.INIT0 = 16'h7888;
    defparam add_4609_27.INIT1 = 16'h7888;
    defparam add_4609_27.INJECT1_0 = "NO";
    defparam add_4609_27.INJECT1_1 = "NO";
    CCU2D add_4609_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[12]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[25]), .B1(nZ0_d2[12]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[13]), .CIN(n61942), .COUT(n61943), .S0(buf_x[1170]), 
          .S1(buf_x[1171]));
    defparam add_4609_25.INIT0 = 16'h7888;
    defparam add_4609_25.INIT1 = 16'h7888;
    defparam add_4609_25.INJECT1_0 = "NO";
    defparam add_4609_25.INJECT1_1 = "NO";
    CCU2D add_4609_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[12]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[23]), .B1(nZ0_d2[12]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[13]), .CIN(n61941), .COUT(n61942), .S0(buf_x[1168]), 
          .S1(buf_x[1169]));
    defparam add_4609_23.INIT0 = 16'h7888;
    defparam add_4609_23.INIT1 = 16'h7888;
    defparam add_4609_23.INJECT1_0 = "NO";
    defparam add_4609_23.INJECT1_1 = "NO";
    CCU2D add_4609_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[12]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[21]), .B1(nZ0_d2[12]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[13]), .CIN(n61940), .COUT(n61941), .S0(buf_x[1166]), 
          .S1(buf_x[1167]));
    defparam add_4609_21.INIT0 = 16'h7888;
    defparam add_4609_21.INIT1 = 16'h7888;
    defparam add_4609_21.INJECT1_0 = "NO";
    defparam add_4609_21.INJECT1_1 = "NO";
    CCU2D add_4609_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[12]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[19]), .B1(nZ0_d2[12]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[13]), .CIN(n61939), .COUT(n61940), .S0(buf_x[1164]), 
          .S1(buf_x[1165]));
    defparam add_4609_19.INIT0 = 16'h7888;
    defparam add_4609_19.INIT1 = 16'h7888;
    defparam add_4609_19.INJECT1_0 = "NO";
    defparam add_4609_19.INJECT1_1 = "NO";
    CCU2D add_4609_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[12]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[17]), .B1(nZ0_d2[12]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[13]), .CIN(n61938), .COUT(n61939), .S0(buf_x[1162]), 
          .S1(buf_x[1163]));
    defparam add_4609_17.INIT0 = 16'h7888;
    defparam add_4609_17.INIT1 = 16'h7888;
    defparam add_4609_17.INJECT1_0 = "NO";
    defparam add_4609_17.INJECT1_1 = "NO";
    CCU2D add_4609_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[12]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[15]), .B1(nZ0_d2[12]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[13]), .CIN(n61937), .COUT(n61938), .S0(buf_x[1160]), 
          .S1(buf_x[1161]));
    defparam add_4609_15.INIT0 = 16'h7888;
    defparam add_4609_15.INIT1 = 16'h7888;
    defparam add_4609_15.INJECT1_0 = "NO";
    defparam add_4609_15.INJECT1_1 = "NO";
    CCU2D add_4609_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[12]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[13]), .B1(nZ0_d2[12]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[13]), .CIN(n61936), .COUT(n61937), .S0(buf_x[1158]), 
          .S1(buf_x[1159]));
    defparam add_4609_13.INIT0 = 16'h7888;
    defparam add_4609_13.INIT1 = 16'h7888;
    defparam add_4609_13.INJECT1_0 = "NO";
    defparam add_4609_13.INJECT1_1 = "NO";
    CCU2D add_4609_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[12]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[11]), .B1(nZ0_d2[12]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[13]), .CIN(n61935), .COUT(n61936), .S0(buf_x[1156]), 
          .S1(buf_x[1157]));
    defparam add_4609_11.INIT0 = 16'h7888;
    defparam add_4609_11.INIT1 = 16'h7888;
    defparam add_4609_11.INJECT1_0 = "NO";
    defparam add_4609_11.INJECT1_1 = "NO";
    CCU2D add_4609_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[12]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[9]), .B1(nZ0_d2[12]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[13]), .CIN(n61934), .COUT(n61935), .S0(buf_x[1154]), 
          .S1(buf_x[1155]));
    defparam add_4609_9.INIT0 = 16'h7888;
    defparam add_4609_9.INIT1 = 16'h7888;
    defparam add_4609_9.INJECT1_0 = "NO";
    defparam add_4609_9.INJECT1_1 = "NO";
    CCU2D add_4609_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[12]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[7]), .B1(nZ0_d2[12]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[13]), .CIN(n61933), .COUT(n61934), .S0(buf_x[1152]), 
          .S1(buf_x[1153]));
    defparam add_4609_7.INIT0 = 16'h7888;
    defparam add_4609_7.INIT1 = 16'h7888;
    defparam add_4609_7.INJECT1_0 = "NO";
    defparam add_4609_7.INJECT1_1 = "NO";
    CCU2D add_4609_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[12]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[5]), .B1(nZ0_d2[12]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[13]), .CIN(n61932), .COUT(n61933), .S0(buf_x[1150]), 
          .S1(buf_x[1151]));
    defparam add_4609_5.INIT0 = 16'h7888;
    defparam add_4609_5.INIT1 = 16'h7888;
    defparam add_4609_5.INJECT1_0 = "NO";
    defparam add_4609_5.INJECT1_1 = "NO";
    CCU2D add_4609_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[12]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[13]), .A1(nEY1_d2[3]), .B1(nZ0_d2[12]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[13]), .CIN(n61931), .COUT(n61932), .S0(buf_x[1148]), 
          .S1(buf_x[1149]));
    defparam add_4609_3.INIT0 = 16'h7888;
    defparam add_4609_3.INIT1 = 16'h7888;
    defparam add_4609_3.INJECT1_0 = "NO";
    defparam add_4609_3.INJECT1_1 = "NO";
    CCU2D add_4609_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[12]), .C1(nEY1_d2[0]), .D1(nZ0_d2[13]), 
          .COUT(n61931), .S1(buf_x[1147]));
    defparam add_4609_1.INIT0 = 16'hF000;
    defparam add_4609_1.INIT1 = 16'h7888;
    defparam add_4609_1.INJECT1_0 = "NO";
    defparam add_4609_1.INJECT1_1 = "NO";
    CCU2D add_4608_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[11]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61930), .S0(buf_x[1143]), .S1(buf_x[1144]));
    defparam add_4608_29.INIT0 = 16'h7888;
    defparam add_4608_29.INIT1 = 16'h0000;
    defparam add_4608_29.INJECT1_0 = "NO";
    defparam add_4608_29.INJECT1_1 = "NO";
    CCU2D add_4608_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[10]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[27]), .B1(nZ0_d2[10]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[11]), .CIN(n61929), .COUT(n61930), .S0(buf_x[1141]), 
          .S1(buf_x[1142]));
    defparam add_4608_27.INIT0 = 16'h7888;
    defparam add_4608_27.INIT1 = 16'h7888;
    defparam add_4608_27.INJECT1_0 = "NO";
    defparam add_4608_27.INJECT1_1 = "NO";
    CCU2D add_4608_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[10]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[25]), .B1(nZ0_d2[10]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[11]), .CIN(n61928), .COUT(n61929), .S0(buf_x[1139]), 
          .S1(buf_x[1140]));
    defparam add_4608_25.INIT0 = 16'h7888;
    defparam add_4608_25.INIT1 = 16'h7888;
    defparam add_4608_25.INJECT1_0 = "NO";
    defparam add_4608_25.INJECT1_1 = "NO";
    CCU2D add_4608_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[10]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[23]), .B1(nZ0_d2[10]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[11]), .CIN(n61927), .COUT(n61928), .S0(buf_x[1137]), 
          .S1(buf_x[1138]));
    defparam add_4608_23.INIT0 = 16'h7888;
    defparam add_4608_23.INIT1 = 16'h7888;
    defparam add_4608_23.INJECT1_0 = "NO";
    defparam add_4608_23.INJECT1_1 = "NO";
    CCU2D add_4608_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[10]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[21]), .B1(nZ0_d2[10]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[11]), .CIN(n61926), .COUT(n61927), .S0(buf_x[1135]), 
          .S1(buf_x[1136]));
    defparam add_4608_21.INIT0 = 16'h7888;
    defparam add_4608_21.INIT1 = 16'h7888;
    defparam add_4608_21.INJECT1_0 = "NO";
    defparam add_4608_21.INJECT1_1 = "NO";
    CCU2D add_4608_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[10]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[19]), .B1(nZ0_d2[10]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[11]), .CIN(n61925), .COUT(n61926), .S0(buf_x[1133]), 
          .S1(buf_x[1134]));
    defparam add_4608_19.INIT0 = 16'h7888;
    defparam add_4608_19.INIT1 = 16'h7888;
    defparam add_4608_19.INJECT1_0 = "NO";
    defparam add_4608_19.INJECT1_1 = "NO";
    CCU2D add_4608_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[10]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[17]), .B1(nZ0_d2[10]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[11]), .CIN(n61924), .COUT(n61925), .S0(buf_x[1131]), 
          .S1(buf_x[1132]));
    defparam add_4608_17.INIT0 = 16'h7888;
    defparam add_4608_17.INIT1 = 16'h7888;
    defparam add_4608_17.INJECT1_0 = "NO";
    defparam add_4608_17.INJECT1_1 = "NO";
    CCU2D add_4608_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[10]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[15]), .B1(nZ0_d2[10]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[11]), .CIN(n61923), .COUT(n61924), .S0(buf_x[1129]), 
          .S1(buf_x[1130]));
    defparam add_4608_15.INIT0 = 16'h7888;
    defparam add_4608_15.INIT1 = 16'h7888;
    defparam add_4608_15.INJECT1_0 = "NO";
    defparam add_4608_15.INJECT1_1 = "NO";
    CCU2D add_4608_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[10]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[13]), .B1(nZ0_d2[10]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[11]), .CIN(n61922), .COUT(n61923), .S0(buf_x[1127]), 
          .S1(buf_x[1128]));
    defparam add_4608_13.INIT0 = 16'h7888;
    defparam add_4608_13.INIT1 = 16'h7888;
    defparam add_4608_13.INJECT1_0 = "NO";
    defparam add_4608_13.INJECT1_1 = "NO";
    CCU2D add_4608_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[10]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[11]), .B1(nZ0_d2[10]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[11]), .CIN(n61921), .COUT(n61922), .S0(buf_x[1125]), 
          .S1(buf_x[1126]));
    defparam add_4608_11.INIT0 = 16'h7888;
    defparam add_4608_11.INIT1 = 16'h7888;
    defparam add_4608_11.INJECT1_0 = "NO";
    defparam add_4608_11.INJECT1_1 = "NO";
    CCU2D add_4608_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[10]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[9]), .B1(nZ0_d2[10]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[11]), .CIN(n61920), .COUT(n61921), .S0(buf_x[1123]), 
          .S1(buf_x[1124]));
    defparam add_4608_9.INIT0 = 16'h7888;
    defparam add_4608_9.INIT1 = 16'h7888;
    defparam add_4608_9.INJECT1_0 = "NO";
    defparam add_4608_9.INJECT1_1 = "NO";
    CCU2D add_4608_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[10]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[7]), .B1(nZ0_d2[10]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[11]), .CIN(n61919), .COUT(n61920), .S0(buf_x[1121]), 
          .S1(buf_x[1122]));
    defparam add_4608_7.INIT0 = 16'h7888;
    defparam add_4608_7.INIT1 = 16'h7888;
    defparam add_4608_7.INJECT1_0 = "NO";
    defparam add_4608_7.INJECT1_1 = "NO";
    CCU2D add_4608_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[10]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[5]), .B1(nZ0_d2[10]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[11]), .CIN(n61918), .COUT(n61919), .S0(buf_x[1119]), 
          .S1(buf_x[1120]));
    defparam add_4608_5.INIT0 = 16'h7888;
    defparam add_4608_5.INIT1 = 16'h7888;
    defparam add_4608_5.INJECT1_0 = "NO";
    defparam add_4608_5.INJECT1_1 = "NO";
    CCU2D add_4608_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[10]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[11]), .A1(nEY1_d2[3]), .B1(nZ0_d2[10]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[11]), .CIN(n61917), .COUT(n61918), .S0(buf_x[1117]), 
          .S1(buf_x[1118]));
    defparam add_4608_3.INIT0 = 16'h7888;
    defparam add_4608_3.INIT1 = 16'h7888;
    defparam add_4608_3.INJECT1_0 = "NO";
    defparam add_4608_3.INJECT1_1 = "NO";
    CCU2D add_4608_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[10]), .C1(nEY1_d2[0]), .D1(nZ0_d2[11]), 
          .COUT(n61917), .S1(buf_x[1116]));
    defparam add_4608_1.INIT0 = 16'hF000;
    defparam add_4608_1.INIT1 = 16'h7888;
    defparam add_4608_1.INJECT1_0 = "NO";
    defparam add_4608_1.INJECT1_1 = "NO";
    CCU2D add_4607_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[9]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61916), .S0(buf_x[1112]), .S1(buf_x[1113]));
    defparam add_4607_29.INIT0 = 16'h7888;
    defparam add_4607_29.INIT1 = 16'h0000;
    defparam add_4607_29.INJECT1_0 = "NO";
    defparam add_4607_29.INJECT1_1 = "NO";
    CCU2D add_4607_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[8]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[27]), .B1(nZ0_d2[8]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[9]), .CIN(n61915), .COUT(n61916), .S0(buf_x[1110]), 
          .S1(buf_x[1111]));
    defparam add_4607_27.INIT0 = 16'h7888;
    defparam add_4607_27.INIT1 = 16'h7888;
    defparam add_4607_27.INJECT1_0 = "NO";
    defparam add_4607_27.INJECT1_1 = "NO";
    CCU2D add_4607_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[8]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[25]), .B1(nZ0_d2[8]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[9]), .CIN(n61914), .COUT(n61915), .S0(buf_x[1108]), 
          .S1(buf_x[1109]));
    defparam add_4607_25.INIT0 = 16'h7888;
    defparam add_4607_25.INIT1 = 16'h7888;
    defparam add_4607_25.INJECT1_0 = "NO";
    defparam add_4607_25.INJECT1_1 = "NO";
    CCU2D add_4607_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[8]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[23]), .B1(nZ0_d2[8]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[9]), .CIN(n61913), .COUT(n61914), .S0(buf_x[1106]), 
          .S1(buf_x[1107]));
    defparam add_4607_23.INIT0 = 16'h7888;
    defparam add_4607_23.INIT1 = 16'h7888;
    defparam add_4607_23.INJECT1_0 = "NO";
    defparam add_4607_23.INJECT1_1 = "NO";
    CCU2D add_4607_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[8]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[21]), .B1(nZ0_d2[8]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[9]), .CIN(n61912), .COUT(n61913), .S0(buf_x[1104]), 
          .S1(buf_x[1105]));
    defparam add_4607_21.INIT0 = 16'h7888;
    defparam add_4607_21.INIT1 = 16'h7888;
    defparam add_4607_21.INJECT1_0 = "NO";
    defparam add_4607_21.INJECT1_1 = "NO";
    CCU2D add_4607_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[8]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[19]), .B1(nZ0_d2[8]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[9]), .CIN(n61911), .COUT(n61912), .S0(buf_x[1102]), 
          .S1(buf_x[1103]));
    defparam add_4607_19.INIT0 = 16'h7888;
    defparam add_4607_19.INIT1 = 16'h7888;
    defparam add_4607_19.INJECT1_0 = "NO";
    defparam add_4607_19.INJECT1_1 = "NO";
    CCU2D add_4607_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[8]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[17]), .B1(nZ0_d2[8]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[9]), .CIN(n61910), .COUT(n61911), .S0(buf_x[1100]), 
          .S1(buf_x[1101]));
    defparam add_4607_17.INIT0 = 16'h7888;
    defparam add_4607_17.INIT1 = 16'h7888;
    defparam add_4607_17.INJECT1_0 = "NO";
    defparam add_4607_17.INJECT1_1 = "NO";
    CCU2D add_4607_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[8]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[15]), .B1(nZ0_d2[8]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[9]), .CIN(n61909), .COUT(n61910), .S0(buf_x[1098]), 
          .S1(buf_x[1099]));
    defparam add_4607_15.INIT0 = 16'h7888;
    defparam add_4607_15.INIT1 = 16'h7888;
    defparam add_4607_15.INJECT1_0 = "NO";
    defparam add_4607_15.INJECT1_1 = "NO";
    CCU2D add_4607_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[8]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[13]), .B1(nZ0_d2[8]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[9]), .CIN(n61908), .COUT(n61909), .S0(buf_x[1096]), 
          .S1(buf_x[1097]));
    defparam add_4607_13.INIT0 = 16'h7888;
    defparam add_4607_13.INIT1 = 16'h7888;
    defparam add_4607_13.INJECT1_0 = "NO";
    defparam add_4607_13.INJECT1_1 = "NO";
    CCU2D add_4607_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[8]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[11]), .B1(nZ0_d2[8]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[9]), .CIN(n61907), .COUT(n61908), .S0(buf_x[1094]), 
          .S1(buf_x[1095]));
    defparam add_4607_11.INIT0 = 16'h7888;
    defparam add_4607_11.INIT1 = 16'h7888;
    defparam add_4607_11.INJECT1_0 = "NO";
    defparam add_4607_11.INJECT1_1 = "NO";
    CCU2D add_4607_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[8]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[9]), .B1(nZ0_d2[8]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[9]), .CIN(n61906), .COUT(n61907), .S0(buf_x[1092]), 
          .S1(buf_x[1093]));
    defparam add_4607_9.INIT0 = 16'h7888;
    defparam add_4607_9.INIT1 = 16'h7888;
    defparam add_4607_9.INJECT1_0 = "NO";
    defparam add_4607_9.INJECT1_1 = "NO";
    CCU2D add_4607_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[8]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[7]), .B1(nZ0_d2[8]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[9]), .CIN(n61905), .COUT(n61906), .S0(buf_x[1090]), 
          .S1(buf_x[1091]));
    defparam add_4607_7.INIT0 = 16'h7888;
    defparam add_4607_7.INIT1 = 16'h7888;
    defparam add_4607_7.INJECT1_0 = "NO";
    defparam add_4607_7.INJECT1_1 = "NO";
    CCU2D add_4607_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[8]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[5]), .B1(nZ0_d2[8]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[9]), .CIN(n61904), .COUT(n61905), .S0(buf_x[1088]), 
          .S1(buf_x[1089]));
    defparam add_4607_5.INIT0 = 16'h7888;
    defparam add_4607_5.INIT1 = 16'h7888;
    defparam add_4607_5.INJECT1_0 = "NO";
    defparam add_4607_5.INJECT1_1 = "NO";
    CCU2D add_4607_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[8]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[9]), .A1(nEY1_d2[3]), .B1(nZ0_d2[8]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[9]), .CIN(n61903), .COUT(n61904), .S0(buf_x[1086]), 
          .S1(buf_x[1087]));
    defparam add_4607_3.INIT0 = 16'h7888;
    defparam add_4607_3.INIT1 = 16'h7888;
    defparam add_4607_3.INJECT1_0 = "NO";
    defparam add_4607_3.INJECT1_1 = "NO";
    CCU2D add_4607_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[8]), .C1(nEY1_d2[0]), .D1(nZ0_d2[9]), 
          .COUT(n61903), .S1(buf_x[1085]));
    defparam add_4607_1.INIT0 = 16'hF000;
    defparam add_4607_1.INIT1 = 16'h7888;
    defparam add_4607_1.INJECT1_0 = "NO";
    defparam add_4607_1.INJECT1_1 = "NO";
    CCU2D add_4606_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[7]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61902), .S0(buf_x[1081]), .S1(buf_x[1082]));
    defparam add_4606_29.INIT0 = 16'h7888;
    defparam add_4606_29.INIT1 = 16'h0000;
    defparam add_4606_29.INJECT1_0 = "NO";
    defparam add_4606_29.INJECT1_1 = "NO";
    CCU2D add_4606_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[6]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[27]), .B1(nZ0_d2[6]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[7]), .CIN(n61901), .COUT(n61902), .S0(buf_x[1079]), 
          .S1(buf_x[1080]));
    defparam add_4606_27.INIT0 = 16'h7888;
    defparam add_4606_27.INIT1 = 16'h7888;
    defparam add_4606_27.INJECT1_0 = "NO";
    defparam add_4606_27.INJECT1_1 = "NO";
    CCU2D add_4606_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[6]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[25]), .B1(nZ0_d2[6]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[7]), .CIN(n61900), .COUT(n61901), .S0(buf_x[1077]), 
          .S1(buf_x[1078]));
    defparam add_4606_25.INIT0 = 16'h7888;
    defparam add_4606_25.INIT1 = 16'h7888;
    defparam add_4606_25.INJECT1_0 = "NO";
    defparam add_4606_25.INJECT1_1 = "NO";
    CCU2D add_4606_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[6]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[23]), .B1(nZ0_d2[6]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[7]), .CIN(n61899), .COUT(n61900), .S0(buf_x[1075]), 
          .S1(buf_x[1076]));
    defparam add_4606_23.INIT0 = 16'h7888;
    defparam add_4606_23.INIT1 = 16'h7888;
    defparam add_4606_23.INJECT1_0 = "NO";
    defparam add_4606_23.INJECT1_1 = "NO";
    CCU2D add_4606_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[6]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[21]), .B1(nZ0_d2[6]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[7]), .CIN(n61898), .COUT(n61899), .S0(buf_x[1073]), 
          .S1(buf_x[1074]));
    defparam add_4606_21.INIT0 = 16'h7888;
    defparam add_4606_21.INIT1 = 16'h7888;
    defparam add_4606_21.INJECT1_0 = "NO";
    defparam add_4606_21.INJECT1_1 = "NO";
    CCU2D add_4606_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[6]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[19]), .B1(nZ0_d2[6]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[7]), .CIN(n61897), .COUT(n61898), .S0(buf_x[1071]), 
          .S1(buf_x[1072]));
    defparam add_4606_19.INIT0 = 16'h7888;
    defparam add_4606_19.INIT1 = 16'h7888;
    defparam add_4606_19.INJECT1_0 = "NO";
    defparam add_4606_19.INJECT1_1 = "NO";
    CCU2D add_4606_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[6]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[17]), .B1(nZ0_d2[6]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[7]), .CIN(n61896), .COUT(n61897), .S0(buf_x[1069]), 
          .S1(buf_x[1070]));
    defparam add_4606_17.INIT0 = 16'h7888;
    defparam add_4606_17.INIT1 = 16'h7888;
    defparam add_4606_17.INJECT1_0 = "NO";
    defparam add_4606_17.INJECT1_1 = "NO";
    CCU2D add_4606_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[6]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[15]), .B1(nZ0_d2[6]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[7]), .CIN(n61895), .COUT(n61896), .S0(buf_x[1067]), 
          .S1(buf_x[1068]));
    defparam add_4606_15.INIT0 = 16'h7888;
    defparam add_4606_15.INIT1 = 16'h7888;
    defparam add_4606_15.INJECT1_0 = "NO";
    defparam add_4606_15.INJECT1_1 = "NO";
    CCU2D add_4606_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[6]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[13]), .B1(nZ0_d2[6]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[7]), .CIN(n61894), .COUT(n61895), .S0(buf_x[1065]), 
          .S1(buf_x[1066]));
    defparam add_4606_13.INIT0 = 16'h7888;
    defparam add_4606_13.INIT1 = 16'h7888;
    defparam add_4606_13.INJECT1_0 = "NO";
    defparam add_4606_13.INJECT1_1 = "NO";
    CCU2D add_4606_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[6]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[11]), .B1(nZ0_d2[6]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[7]), .CIN(n61893), .COUT(n61894), .S0(buf_x[1063]), 
          .S1(buf_x[1064]));
    defparam add_4606_11.INIT0 = 16'h7888;
    defparam add_4606_11.INIT1 = 16'h7888;
    defparam add_4606_11.INJECT1_0 = "NO";
    defparam add_4606_11.INJECT1_1 = "NO";
    CCU2D add_4606_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[6]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[9]), .B1(nZ0_d2[6]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[7]), .CIN(n61892), .COUT(n61893), .S0(buf_x[1061]), 
          .S1(buf_x[1062]));
    defparam add_4606_9.INIT0 = 16'h7888;
    defparam add_4606_9.INIT1 = 16'h7888;
    defparam add_4606_9.INJECT1_0 = "NO";
    defparam add_4606_9.INJECT1_1 = "NO";
    CCU2D add_4606_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[6]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[7]), .B1(nZ0_d2[6]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[7]), .CIN(n61891), .COUT(n61892), .S0(buf_x[1059]), 
          .S1(buf_x[1060]));
    defparam add_4606_7.INIT0 = 16'h7888;
    defparam add_4606_7.INIT1 = 16'h7888;
    defparam add_4606_7.INJECT1_0 = "NO";
    defparam add_4606_7.INJECT1_1 = "NO";
    LUT4 i49853_2_lut (.A(buf_r[1086]), .B(buf_r[1115]), .Z(buf_x[1759])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49853_2_lut.init = 16'h6666;
    CCU2D add_4606_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[6]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[5]), .B1(nZ0_d2[6]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[7]), .CIN(n61890), .COUT(n61891), .S0(buf_x[1057]), 
          .S1(buf_x[1058]));
    defparam add_4606_5.INIT0 = 16'h7888;
    defparam add_4606_5.INIT1 = 16'h7888;
    defparam add_4606_5.INJECT1_0 = "NO";
    defparam add_4606_5.INJECT1_1 = "NO";
    LUT4 i49856_2_lut (.A(buf_x[1526]), .B(buf_x[1555]), .Z(buf_x[1761])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49856_2_lut.init = 16'h6666;
    CCU2D add_4606_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[6]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[7]), .A1(nEY1_d2[3]), .B1(nZ0_d2[6]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[7]), .CIN(n61889), .COUT(n61890), .S0(buf_x[1055]), 
          .S1(buf_x[1056]));
    defparam add_4606_3.INIT0 = 16'h7888;
    defparam add_4606_3.INIT1 = 16'h7888;
    defparam add_4606_3.INJECT1_0 = "NO";
    defparam add_4606_3.INJECT1_1 = "NO";
    LUT4 i49855_2_lut (.A(buf_r[1210]), .B(buf_r[1239]), .Z(buf_x[1796])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49855_2_lut.init = 16'h6666;
    LUT4 i49851_2_lut (.A(buf_x[1592]), .B(buf_x[1621]), .Z(buf_x[1798])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49851_2_lut.init = 16'h6666;
    CCU2D add_4606_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[6]), .C1(nEY1_d2[0]), .D1(nZ0_d2[7]), 
          .COUT(n61889), .S1(buf_x[1054]));
    defparam add_4606_1.INIT0 = 16'hF000;
    defparam add_4606_1.INIT1 = 16'h7888;
    defparam add_4606_1.INJECT1_0 = "NO";
    defparam add_4606_1.INJECT1_1 = "NO";
    CCU2D add_4605_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[5]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61888), .S0(buf_x[1050]), .S1(buf_x[1051]));
    defparam add_4605_29.INIT0 = 16'h7888;
    defparam add_4605_29.INIT1 = 16'h0000;
    defparam add_4605_29.INJECT1_0 = "NO";
    defparam add_4605_29.INJECT1_1 = "NO";
    CCU2D add_4605_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[4]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[27]), .B1(nZ0_d2[4]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[5]), .CIN(n61887), .COUT(n61888), .S0(buf_x[1048]), 
          .S1(buf_x[1049]));
    defparam add_4605_27.INIT0 = 16'h7888;
    defparam add_4605_27.INIT1 = 16'h7888;
    defparam add_4605_27.INJECT1_0 = "NO";
    defparam add_4605_27.INJECT1_1 = "NO";
    CCU2D add_4605_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[4]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[25]), .B1(nZ0_d2[4]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[5]), .CIN(n61886), .COUT(n61887), .S0(buf_x[1046]), 
          .S1(buf_x[1047]));
    defparam add_4605_25.INIT0 = 16'h7888;
    defparam add_4605_25.INIT1 = 16'h7888;
    defparam add_4605_25.INJECT1_0 = "NO";
    defparam add_4605_25.INJECT1_1 = "NO";
    CCU2D add_4605_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[4]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[23]), .B1(nZ0_d2[4]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[5]), .CIN(n61885), .COUT(n61886), .S0(buf_x[1044]), 
          .S1(buf_x[1045]));
    defparam add_4605_23.INIT0 = 16'h7888;
    defparam add_4605_23.INIT1 = 16'h7888;
    defparam add_4605_23.INJECT1_0 = "NO";
    defparam add_4605_23.INJECT1_1 = "NO";
    CCU2D add_4605_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[4]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[21]), .B1(nZ0_d2[4]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[5]), .CIN(n61884), .COUT(n61885), .S0(buf_x[1042]), 
          .S1(buf_x[1043]));
    defparam add_4605_21.INIT0 = 16'h7888;
    defparam add_4605_21.INIT1 = 16'h7888;
    defparam add_4605_21.INJECT1_0 = "NO";
    defparam add_4605_21.INJECT1_1 = "NO";
    CCU2D add_4605_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[4]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[19]), .B1(nZ0_d2[4]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[5]), .CIN(n61883), .COUT(n61884), .S0(buf_x[1040]), 
          .S1(buf_x[1041]));
    defparam add_4605_19.INIT0 = 16'h7888;
    defparam add_4605_19.INIT1 = 16'h7888;
    defparam add_4605_19.INJECT1_0 = "NO";
    defparam add_4605_19.INJECT1_1 = "NO";
    CCU2D add_4605_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[4]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[17]), .B1(nZ0_d2[4]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[5]), .CIN(n61882), .COUT(n61883), .S0(buf_x[1038]), 
          .S1(buf_x[1039]));
    defparam add_4605_17.INIT0 = 16'h7888;
    defparam add_4605_17.INIT1 = 16'h7888;
    defparam add_4605_17.INJECT1_0 = "NO";
    defparam add_4605_17.INJECT1_1 = "NO";
    CCU2D add_4605_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[4]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[15]), .B1(nZ0_d2[4]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[5]), .CIN(n61881), .COUT(n61882), .S0(buf_x[1036]), 
          .S1(buf_x[1037]));
    defparam add_4605_15.INIT0 = 16'h7888;
    defparam add_4605_15.INIT1 = 16'h7888;
    defparam add_4605_15.INJECT1_0 = "NO";
    defparam add_4605_15.INJECT1_1 = "NO";
    CCU2D add_4605_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[4]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[13]), .B1(nZ0_d2[4]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[5]), .CIN(n61880), .COUT(n61881), .S0(buf_x[1034]), 
          .S1(buf_x[1035]));
    defparam add_4605_13.INIT0 = 16'h7888;
    defparam add_4605_13.INIT1 = 16'h7888;
    defparam add_4605_13.INJECT1_0 = "NO";
    defparam add_4605_13.INJECT1_1 = "NO";
    CCU2D add_4605_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[4]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[11]), .B1(nZ0_d2[4]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[5]), .CIN(n61879), .COUT(n61880), .S0(buf_x[1032]), 
          .S1(buf_x[1033]));
    defparam add_4605_11.INIT0 = 16'h7888;
    defparam add_4605_11.INIT1 = 16'h7888;
    defparam add_4605_11.INJECT1_0 = "NO";
    defparam add_4605_11.INJECT1_1 = "NO";
    CCU2D add_4605_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[4]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[9]), .B1(nZ0_d2[4]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[5]), .CIN(n61878), .COUT(n61879), .S0(buf_x[1030]), 
          .S1(buf_x[1031]));
    defparam add_4605_9.INIT0 = 16'h7888;
    defparam add_4605_9.INIT1 = 16'h7888;
    defparam add_4605_9.INJECT1_0 = "NO";
    defparam add_4605_9.INJECT1_1 = "NO";
    CCU2D add_4605_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[4]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[7]), .B1(nZ0_d2[4]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[5]), .CIN(n61877), .COUT(n61878), .S0(buf_x[1028]), 
          .S1(buf_x[1029]));
    defparam add_4605_7.INIT0 = 16'h7888;
    defparam add_4605_7.INIT1 = 16'h7888;
    defparam add_4605_7.INJECT1_0 = "NO";
    defparam add_4605_7.INJECT1_1 = "NO";
    CCU2D add_4605_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[4]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[5]), .B1(nZ0_d2[4]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[5]), .CIN(n61876), .COUT(n61877), .S0(buf_x[1026]), 
          .S1(buf_x[1027]));
    defparam add_4605_5.INIT0 = 16'h7888;
    defparam add_4605_5.INIT1 = 16'h7888;
    defparam add_4605_5.INJECT1_0 = "NO";
    defparam add_4605_5.INJECT1_1 = "NO";
    CCU2D add_4605_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[4]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[5]), .A1(nEY1_d2[3]), .B1(nZ0_d2[4]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[5]), .CIN(n61875), .COUT(n61876), .S0(buf_x[1024]), 
          .S1(buf_x[1025]));
    defparam add_4605_3.INIT0 = 16'h7888;
    defparam add_4605_3.INIT1 = 16'h7888;
    defparam add_4605_3.INJECT1_0 = "NO";
    defparam add_4605_3.INJECT1_1 = "NO";
    CCU2D add_4605_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[4]), .C1(nEY1_d2[0]), .D1(nZ0_d2[5]), 
          .COUT(n61875), .S1(buf_x[1023]));
    defparam add_4605_1.INIT0 = 16'hF000;
    defparam add_4605_1.INIT1 = 16'h7888;
    defparam add_4605_1.INJECT1_0 = "NO";
    defparam add_4605_1.INJECT1_1 = "NO";
    CCU2D add_4604_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[3]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61874), .S0(buf_x[1019]), .S1(buf_x[1020]));
    defparam add_4604_29.INIT0 = 16'h7888;
    defparam add_4604_29.INIT1 = 16'h0000;
    defparam add_4604_29.INJECT1_0 = "NO";
    defparam add_4604_29.INJECT1_1 = "NO";
    CCU2D add_4604_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[2]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[27]), .B1(nZ0_d2[2]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[3]), .CIN(n61873), .COUT(n61874), .S0(buf_x[1017]), 
          .S1(buf_x[1018]));
    defparam add_4604_27.INIT0 = 16'h7888;
    defparam add_4604_27.INIT1 = 16'h7888;
    defparam add_4604_27.INJECT1_0 = "NO";
    defparam add_4604_27.INJECT1_1 = "NO";
    CCU2D add_4604_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[2]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[25]), .B1(nZ0_d2[2]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[3]), .CIN(n61872), .COUT(n61873), .S0(buf_x[1015]), 
          .S1(buf_x[1016]));
    defparam add_4604_25.INIT0 = 16'h7888;
    defparam add_4604_25.INIT1 = 16'h7888;
    defparam add_4604_25.INJECT1_0 = "NO";
    defparam add_4604_25.INJECT1_1 = "NO";
    CCU2D add_4604_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[2]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[23]), .B1(nZ0_d2[2]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[3]), .CIN(n61871), .COUT(n61872), .S0(buf_x[1013]), 
          .S1(buf_x[1014]));
    defparam add_4604_23.INIT0 = 16'h7888;
    defparam add_4604_23.INIT1 = 16'h7888;
    defparam add_4604_23.INJECT1_0 = "NO";
    defparam add_4604_23.INJECT1_1 = "NO";
    CCU2D add_4604_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[2]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[21]), .B1(nZ0_d2[2]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[3]), .CIN(n61870), .COUT(n61871), .S0(buf_x[1011]), 
          .S1(buf_x[1012]));
    defparam add_4604_21.INIT0 = 16'h7888;
    defparam add_4604_21.INIT1 = 16'h7888;
    defparam add_4604_21.INJECT1_0 = "NO";
    defparam add_4604_21.INJECT1_1 = "NO";
    CCU2D add_4604_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[2]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[19]), .B1(nZ0_d2[2]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[3]), .CIN(n61869), .COUT(n61870), .S0(buf_x[1009]), 
          .S1(buf_x[1010]));
    defparam add_4604_19.INIT0 = 16'h7888;
    defparam add_4604_19.INIT1 = 16'h7888;
    defparam add_4604_19.INJECT1_0 = "NO";
    defparam add_4604_19.INJECT1_1 = "NO";
    CCU2D add_4604_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[2]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[17]), .B1(nZ0_d2[2]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[3]), .CIN(n61868), .COUT(n61869), .S0(buf_x[1007]), 
          .S1(buf_x[1008]));
    defparam add_4604_17.INIT0 = 16'h7888;
    defparam add_4604_17.INIT1 = 16'h7888;
    defparam add_4604_17.INJECT1_0 = "NO";
    defparam add_4604_17.INJECT1_1 = "NO";
    CCU2D add_4604_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[2]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[15]), .B1(nZ0_d2[2]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[3]), .CIN(n61867), .COUT(n61868), .S0(buf_x[1005]), 
          .S1(buf_x[1006]));
    defparam add_4604_15.INIT0 = 16'h7888;
    defparam add_4604_15.INIT1 = 16'h7888;
    defparam add_4604_15.INJECT1_0 = "NO";
    defparam add_4604_15.INJECT1_1 = "NO";
    CCU2D add_4604_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[2]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[13]), .B1(nZ0_d2[2]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[3]), .CIN(n61866), .COUT(n61867), .S0(buf_x[1003]), 
          .S1(buf_x[1004]));
    defparam add_4604_13.INIT0 = 16'h7888;
    defparam add_4604_13.INIT1 = 16'h7888;
    defparam add_4604_13.INJECT1_0 = "NO";
    defparam add_4604_13.INJECT1_1 = "NO";
    CCU2D add_4604_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[2]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[11]), .B1(nZ0_d2[2]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[3]), .CIN(n61865), .COUT(n61866), .S0(buf_x[1001]), 
          .S1(buf_x[1002]));
    defparam add_4604_11.INIT0 = 16'h7888;
    defparam add_4604_11.INIT1 = 16'h7888;
    defparam add_4604_11.INJECT1_0 = "NO";
    defparam add_4604_11.INJECT1_1 = "NO";
    CCU2D add_4604_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[2]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[9]), .B1(nZ0_d2[2]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[3]), .CIN(n61864), .COUT(n61865), .S0(buf_x[999]), 
          .S1(buf_x[1000]));
    defparam add_4604_9.INIT0 = 16'h7888;
    defparam add_4604_9.INIT1 = 16'h7888;
    defparam add_4604_9.INJECT1_0 = "NO";
    defparam add_4604_9.INJECT1_1 = "NO";
    CCU2D add_4604_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[2]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[7]), .B1(nZ0_d2[2]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[3]), .CIN(n61863), .COUT(n61864), .S0(buf_x[997]), 
          .S1(buf_x[998]));
    defparam add_4604_7.INIT0 = 16'h7888;
    defparam add_4604_7.INIT1 = 16'h7888;
    defparam add_4604_7.INJECT1_0 = "NO";
    defparam add_4604_7.INJECT1_1 = "NO";
    CCU2D add_4604_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[2]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[5]), .B1(nZ0_d2[2]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[3]), .CIN(n61862), .COUT(n61863), .S0(buf_x[995]), 
          .S1(buf_x[996]));
    defparam add_4604_5.INIT0 = 16'h7888;
    defparam add_4604_5.INIT1 = 16'h7888;
    defparam add_4604_5.INJECT1_0 = "NO";
    defparam add_4604_5.INJECT1_1 = "NO";
    CCU2D add_4604_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[2]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[3]), .A1(nEY1_d2[3]), .B1(nZ0_d2[2]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[3]), .CIN(n61861), .COUT(n61862), .S0(buf_x[993]), 
          .S1(buf_x[994]));
    defparam add_4604_3.INIT0 = 16'h7888;
    defparam add_4604_3.INIT1 = 16'h7888;
    defparam add_4604_3.INJECT1_0 = "NO";
    defparam add_4604_3.INJECT1_1 = "NO";
    CCU2D add_4604_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[2]), .C1(nEY1_d2[0]), .D1(nZ0_d2[3]), 
          .COUT(n61861), .S1(buf_x[992]));
    defparam add_4604_1.INIT0 = 16'hF000;
    defparam add_4604_1.INIT1 = 16'h7888;
    defparam add_4604_1.INJECT1_0 = "NO";
    defparam add_4604_1.INJECT1_1 = "NO";
    CCU2D add_2957_30 (.A0(buf_x[1620]), .B0(buf_x[1649]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1620]), .B1(buf_x[1650]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61854), .S0(buf_x[1826]), .S1(buf_x[1827]));
    defparam add_2957_30.INIT0 = 16'h5666;
    defparam add_2957_30.INIT1 = 16'h5666;
    defparam add_2957_30.INJECT1_0 = "NO";
    defparam add_2957_30.INJECT1_1 = "NO";
    CCU2D add_2957_28 (.A0(buf_x[1618]), .B0(buf_x[1647]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1619]), .B1(buf_x[1648]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61853), .COUT(n61854), .S0(buf_x[1824]), 
          .S1(buf_x[1825]));
    defparam add_2957_28.INIT0 = 16'h5666;
    defparam add_2957_28.INIT1 = 16'h5666;
    defparam add_2957_28.INJECT1_0 = "NO";
    defparam add_2957_28.INJECT1_1 = "NO";
    CCU2D add_2957_26 (.A0(buf_x[1616]), .B0(buf_x[1645]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1617]), .B1(buf_x[1646]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61852), .COUT(n61853), .S0(buf_x[1822]), 
          .S1(buf_x[1823]));
    defparam add_2957_26.INIT0 = 16'h5666;
    defparam add_2957_26.INIT1 = 16'h5666;
    defparam add_2957_26.INJECT1_0 = "NO";
    defparam add_2957_26.INJECT1_1 = "NO";
    CCU2D add_2957_24 (.A0(buf_x[1614]), .B0(buf_x[1643]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1615]), .B1(buf_x[1644]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61851), .COUT(n61852), .S0(buf_x[1820]), 
          .S1(buf_x[1821]));
    defparam add_2957_24.INIT0 = 16'h5666;
    defparam add_2957_24.INIT1 = 16'h5666;
    defparam add_2957_24.INJECT1_0 = "NO";
    defparam add_2957_24.INJECT1_1 = "NO";
    CCU2D add_2957_22 (.A0(buf_x[1612]), .B0(buf_x[1641]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1613]), .B1(buf_x[1642]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61850), .COUT(n61851), .S0(buf_x[1818]), 
          .S1(buf_x[1819]));
    defparam add_2957_22.INIT0 = 16'h5666;
    defparam add_2957_22.INIT1 = 16'h5666;
    defparam add_2957_22.INJECT1_0 = "NO";
    defparam add_2957_22.INJECT1_1 = "NO";
    CCU2D add_2957_20 (.A0(buf_x[1610]), .B0(buf_x[1639]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1611]), .B1(buf_x[1640]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61849), .COUT(n61850), .S0(buf_x[1816]), 
          .S1(buf_x[1817]));
    defparam add_2957_20.INIT0 = 16'h5666;
    defparam add_2957_20.INIT1 = 16'h5666;
    defparam add_2957_20.INJECT1_0 = "NO";
    defparam add_2957_20.INJECT1_1 = "NO";
    CCU2D add_2957_18 (.A0(buf_x[1608]), .B0(buf_x[1637]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1609]), .B1(buf_x[1638]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61848), .COUT(n61849), .S0(buf_x[1814]), 
          .S1(buf_x[1815]));
    defparam add_2957_18.INIT0 = 16'h5666;
    defparam add_2957_18.INIT1 = 16'h5666;
    defparam add_2957_18.INJECT1_0 = "NO";
    defparam add_2957_18.INJECT1_1 = "NO";
    CCU2D add_2957_16 (.A0(buf_x[1606]), .B0(buf_x[1635]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1607]), .B1(buf_x[1636]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61847), .COUT(n61848), .S0(buf_x[1812]), 
          .S1(buf_x[1813]));
    defparam add_2957_16.INIT0 = 16'h5666;
    defparam add_2957_16.INIT1 = 16'h5666;
    defparam add_2957_16.INJECT1_0 = "NO";
    defparam add_2957_16.INJECT1_1 = "NO";
    CCU2D add_2957_14 (.A0(buf_x[1604]), .B0(buf_x[1633]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1605]), .B1(buf_x[1634]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61846), .COUT(n61847), .S0(buf_x[1810]), 
          .S1(buf_x[1811]));
    defparam add_2957_14.INIT0 = 16'h5666;
    defparam add_2957_14.INIT1 = 16'h5666;
    defparam add_2957_14.INJECT1_0 = "NO";
    defparam add_2957_14.INJECT1_1 = "NO";
    CCU2D add_2957_12 (.A0(buf_x[1602]), .B0(buf_x[1631]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1603]), .B1(buf_x[1632]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61845), .COUT(n61846), .S0(buf_x[1808]), 
          .S1(buf_x[1809]));
    defparam add_2957_12.INIT0 = 16'h5666;
    defparam add_2957_12.INIT1 = 16'h5666;
    defparam add_2957_12.INJECT1_0 = "NO";
    defparam add_2957_12.INJECT1_1 = "NO";
    CCU2D add_2957_10 (.A0(buf_x[1600]), .B0(buf_x[1629]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1601]), .B1(buf_x[1630]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61844), .COUT(n61845), .S0(buf_x[1806]), 
          .S1(buf_x[1807]));
    defparam add_2957_10.INIT0 = 16'h5666;
    defparam add_2957_10.INIT1 = 16'h5666;
    defparam add_2957_10.INJECT1_0 = "NO";
    defparam add_2957_10.INJECT1_1 = "NO";
    CCU2D add_2957_8 (.A0(buf_x[1598]), .B0(buf_x[1627]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1599]), .B1(buf_x[1628]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61843), .COUT(n61844), .S0(buf_x[1804]), 
          .S1(buf_x[1805]));
    defparam add_2957_8.INIT0 = 16'h5666;
    defparam add_2957_8.INIT1 = 16'h5666;
    defparam add_2957_8.INJECT1_0 = "NO";
    defparam add_2957_8.INJECT1_1 = "NO";
    CCU2D add_2957_6 (.A0(buf_x[1596]), .B0(buf_x[1625]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1597]), .B1(buf_x[1626]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61842), .COUT(n61843), .S0(buf_x[1802]), 
          .S1(buf_x[1803]));
    defparam add_2957_6.INIT0 = 16'h5666;
    defparam add_2957_6.INIT1 = 16'h5666;
    defparam add_2957_6.INJECT1_0 = "NO";
    defparam add_2957_6.INJECT1_1 = "NO";
    CCU2D add_2957_4 (.A0(buf_x[1594]), .B0(buf_x[1623]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1595]), .B1(buf_x[1624]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61841), .COUT(n61842), .S0(buf_x[1800]), 
          .S1(buf_x[1801]));
    defparam add_2957_4.INIT0 = 16'h5666;
    defparam add_2957_4.INIT1 = 16'h5666;
    defparam add_2957_4.INJECT1_0 = "NO";
    defparam add_2957_4.INJECT1_1 = "NO";
    CCU2D add_2957_2 (.A0(buf_x[1592]), .B0(buf_x[1621]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1593]), .B1(buf_x[1622]), .C1(GND_net), 
          .D1(GND_net), .COUT(n61841), .S1(buf_x[1799]));
    defparam add_2957_2.INIT0 = 16'h7000;
    defparam add_2957_2.INIT1 = 16'h5666;
    defparam add_2957_2.INJECT1_0 = "NO";
    defparam add_2957_2.INJECT1_1 = "NO";
    FD1S3IX buf_r_991__808 (.D(nEY1_d2[0]), .CK(clock), .CD(n23965), .Q(buf_r[991]));
    defparam buf_r_991__808.GSR = "DISABLED";
    FD1S3IX buf_r_1022__777 (.D(nEY1_d2[0]), .CK(clock), .CD(n23964), 
            .Q(buf_x[1489]));
    defparam buf_r_1022__777.GSR = "DISABLED";
    FD1S3IX buf_r_1053__746 (.D(nEY1_d2[0]), .CK(clock), .CD(n23963), 
            .Q(buf_r[1053]));
    defparam buf_r_1053__746.GSR = "DISABLED";
    FD1S3IX buf_r_1084__715 (.D(nEY1_d2[0]), .CK(clock), .CD(n23962), 
            .Q(buf_x[1757]));
    defparam buf_r_1084__715.GSR = "DISABLED";
    FD1S3IX buf_r_1115__684 (.D(nEY1_d2[0]), .CK(clock), .CD(n23961), 
            .Q(buf_r[1115]));
    defparam buf_r_1115__684.GSR = "DISABLED";
    FD1S3IX buf_r_1146__653 (.D(nEY1_d2[0]), .CK(clock), .CD(n23960), 
            .Q(buf_x[1555]));
    defparam buf_r_1146__653.GSR = "DISABLED";
    FD1S3IX buf_r_1177__622 (.D(nEY1_d2[0]), .CK(clock), .CD(n23959), 
            .Q(buf_r[1177]));
    defparam buf_r_1177__622.GSR = "DISABLED";
    FD1S3IX buf_r_1208__591 (.D(nEY1_d2[0]), .CK(clock), .CD(n23958), 
            .Q(buf_x[1794]));
    defparam buf_r_1208__591.GSR = "DISABLED";
    FD1S3IX buf_r_1239__560 (.D(nEY1_d2[0]), .CK(clock), .CD(n23957), 
            .Q(buf_r[1239]));
    defparam buf_r_1239__560.GSR = "DISABLED";
    FD1S3IX buf_r_1270__529 (.D(nEY1_d2[0]), .CK(clock), .CD(n23956), 
            .Q(buf_x[1621]));
    defparam buf_r_1270__529.GSR = "DISABLED";
    CCU2D add_4603_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[1]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61779), .S0(buf_x[988]), .S1(buf_x[989]));
    defparam add_4603_29.INIT0 = 16'h7888;
    defparam add_4603_29.INIT1 = 16'h0000;
    defparam add_4603_29.INJECT1_0 = "NO";
    defparam add_4603_29.INJECT1_1 = "NO";
    CCU2D add_4603_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[0]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[27]), .B1(nZ0_d2[0]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[1]), .CIN(n61778), .COUT(n61779), .S0(buf_x[986]), 
          .S1(buf_x[987]));
    defparam add_4603_27.INIT0 = 16'h7888;
    defparam add_4603_27.INIT1 = 16'h7888;
    defparam add_4603_27.INJECT1_0 = "NO";
    defparam add_4603_27.INJECT1_1 = "NO";
    CCU2D add_4603_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[0]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[25]), .B1(nZ0_d2[0]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[1]), .CIN(n61777), .COUT(n61778), .S0(buf_x[984]), 
          .S1(buf_x[985]));
    defparam add_4603_25.INIT0 = 16'h7888;
    defparam add_4603_25.INIT1 = 16'h7888;
    defparam add_4603_25.INJECT1_0 = "NO";
    defparam add_4603_25.INJECT1_1 = "NO";
    CCU2D add_4603_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[0]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[23]), .B1(nZ0_d2[0]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[1]), .CIN(n61776), .COUT(n61777), .S0(buf_x[982]), 
          .S1(buf_x[983]));
    defparam add_4603_23.INIT0 = 16'h7888;
    defparam add_4603_23.INIT1 = 16'h7888;
    defparam add_4603_23.INJECT1_0 = "NO";
    defparam add_4603_23.INJECT1_1 = "NO";
    CCU2D add_4603_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[0]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[21]), .B1(nZ0_d2[0]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[1]), .CIN(n61775), .COUT(n61776), .S0(buf_x[980]), 
          .S1(buf_x[981]));
    defparam add_4603_21.INIT0 = 16'h7888;
    defparam add_4603_21.INIT1 = 16'h7888;
    defparam add_4603_21.INJECT1_0 = "NO";
    defparam add_4603_21.INJECT1_1 = "NO";
    CCU2D add_4603_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[0]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[19]), .B1(nZ0_d2[0]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[1]), .CIN(n61774), .COUT(n61775), .S0(buf_x[978]), 
          .S1(buf_x[979]));
    defparam add_4603_19.INIT0 = 16'h7888;
    defparam add_4603_19.INIT1 = 16'h7888;
    defparam add_4603_19.INJECT1_0 = "NO";
    defparam add_4603_19.INJECT1_1 = "NO";
    CCU2D add_4603_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[0]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[17]), .B1(nZ0_d2[0]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[1]), .CIN(n61773), .COUT(n61774), .S0(buf_x[976]), 
          .S1(buf_x[977]));
    defparam add_4603_17.INIT0 = 16'h7888;
    defparam add_4603_17.INIT1 = 16'h7888;
    defparam add_4603_17.INJECT1_0 = "NO";
    defparam add_4603_17.INJECT1_1 = "NO";
    CCU2D add_4603_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[0]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[15]), .B1(nZ0_d2[0]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[1]), .CIN(n61772), .COUT(n61773), .S0(buf_x[974]), 
          .S1(buf_x[975]));
    defparam add_4603_15.INIT0 = 16'h7888;
    defparam add_4603_15.INIT1 = 16'h7888;
    defparam add_4603_15.INJECT1_0 = "NO";
    defparam add_4603_15.INJECT1_1 = "NO";
    CCU2D add_4603_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[0]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[13]), .B1(nZ0_d2[0]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[1]), .CIN(n61771), .COUT(n61772), .S0(buf_x[972]), 
          .S1(buf_x[973]));
    defparam add_4603_13.INIT0 = 16'h7888;
    defparam add_4603_13.INIT1 = 16'h7888;
    defparam add_4603_13.INJECT1_0 = "NO";
    defparam add_4603_13.INJECT1_1 = "NO";
    CCU2D add_4603_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[0]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[11]), .B1(nZ0_d2[0]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[1]), .CIN(n61770), .COUT(n61771), .S0(buf_x[970]), 
          .S1(buf_x[971]));
    defparam add_4603_11.INIT0 = 16'h7888;
    defparam add_4603_11.INIT1 = 16'h7888;
    defparam add_4603_11.INJECT1_0 = "NO";
    defparam add_4603_11.INJECT1_1 = "NO";
    CCU2D add_4603_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[0]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[9]), .B1(nZ0_d2[0]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[1]), .CIN(n61769), .COUT(n61770), .S0(buf_x[968]), 
          .S1(buf_x[969]));
    defparam add_4603_9.INIT0 = 16'h7888;
    defparam add_4603_9.INIT1 = 16'h7888;
    defparam add_4603_9.INJECT1_0 = "NO";
    defparam add_4603_9.INJECT1_1 = "NO";
    CCU2D add_4603_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[0]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[7]), .B1(nZ0_d2[0]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[1]), .CIN(n61768), .COUT(n61769), .S0(buf_x[966]), 
          .S1(buf_x[967]));
    defparam add_4603_7.INIT0 = 16'h7888;
    defparam add_4603_7.INIT1 = 16'h7888;
    defparam add_4603_7.INJECT1_0 = "NO";
    defparam add_4603_7.INJECT1_1 = "NO";
    CCU2D add_4603_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[0]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[5]), .B1(nZ0_d2[0]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[1]), .CIN(n61767), .COUT(n61768), .S0(buf_x[964]), 
          .S1(buf_x[965]));
    defparam add_4603_5.INIT0 = 16'h7888;
    defparam add_4603_5.INIT1 = 16'h7888;
    defparam add_4603_5.INJECT1_0 = "NO";
    defparam add_4603_5.INJECT1_1 = "NO";
    CCU2D add_4603_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[0]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[1]), .A1(nEY1_d2[3]), .B1(nZ0_d2[0]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[1]), .CIN(n61766), .COUT(n61767), .S0(buf_x[962]), 
          .S1(buf_x[963]));
    defparam add_4603_3.INIT0 = 16'h7888;
    defparam add_4603_3.INIT1 = 16'h7888;
    defparam add_4603_3.INJECT1_0 = "NO";
    defparam add_4603_3.INJECT1_1 = "NO";
    CCU2D add_4603_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[0]), .C1(nEY1_d2[0]), .D1(nZ0_d2[1]), 
          .COUT(n61766));
    defparam add_4603_1.INIT0 = 16'hF000;
    defparam add_4603_1.INIT1 = 16'h7888;
    defparam add_4603_1.INJECT1_0 = "NO";
    defparam add_4603_1.INJECT1_1 = "NO";
    CCU2D add_952_34 (.A0(buf_x[1912]), .B0(buf_x[1945]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1912]), .B1(buf_x[1946]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62154), .S0(\nZ1_e0[48] ), .S1(\nZ1_e0[49] ));
    defparam add_952_34.INIT0 = 16'h5666;
    defparam add_952_34.INIT1 = 16'h5666;
    defparam add_952_34.INJECT1_0 = "NO";
    defparam add_952_34.INJECT1_1 = "NO";
    CCU2D add_952_32 (.A0(buf_x[1912]), .B0(buf_x[1943]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1912]), .B1(buf_x[1944]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62153), .COUT(n62154), .S0(\nZ1_e0[46] ), 
          .S1(\nZ1_e0[47] ));
    defparam add_952_32.INIT0 = 16'h5666;
    defparam add_952_32.INIT1 = 16'h5666;
    defparam add_952_32.INJECT1_0 = "NO";
    defparam add_952_32.INJECT1_1 = "NO";
    CCU2D add_952_30 (.A0(buf_x[1912]), .B0(buf_x[1941]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1912]), .B1(buf_x[1942]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62152), .COUT(n62153), .S0(\nZ1_e0[44] ), 
          .S1(\nZ1_e0[45] ));
    defparam add_952_30.INIT0 = 16'h5666;
    defparam add_952_30.INIT1 = 16'h5666;
    defparam add_952_30.INJECT1_0 = "NO";
    defparam add_952_30.INJECT1_1 = "NO";
    CCU2D add_952_28 (.A0(buf_x[1910]), .B0(buf_x[1939]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1911]), .B1(buf_x[1940]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62151), .COUT(n62152), .S0(\nZ1_e0[42] ), 
          .S1(\nZ1_e0[43] ));
    defparam add_952_28.INIT0 = 16'h5666;
    defparam add_952_28.INIT1 = 16'h5666;
    defparam add_952_28.INJECT1_0 = "NO";
    defparam add_952_28.INJECT1_1 = "NO";
    CCU2D add_952_26 (.A0(buf_x[1908]), .B0(buf_x[1937]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1909]), .B1(buf_x[1938]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62150), .COUT(n62151), .S0(\nZ1_e0[40] ), 
          .S1(\nZ1_e0[41] ));
    defparam add_952_26.INIT0 = 16'h5666;
    defparam add_952_26.INIT1 = 16'h5666;
    defparam add_952_26.INJECT1_0 = "NO";
    defparam add_952_26.INJECT1_1 = "NO";
    CCU2D add_952_24 (.A0(buf_x[1906]), .B0(buf_x[1935]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1907]), .B1(buf_x[1936]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62149), .COUT(n62150), .S0(\nZ1_e0[38] ), 
          .S1(\nZ1_e0[39] ));
    defparam add_952_24.INIT0 = 16'h5666;
    defparam add_952_24.INIT1 = 16'h5666;
    defparam add_952_24.INJECT1_0 = "NO";
    defparam add_952_24.INJECT1_1 = "NO";
    CCU2D add_952_22 (.A0(buf_x[1904]), .B0(buf_x[1933]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1905]), .B1(buf_x[1934]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62148), .COUT(n62149), .S0(\nZ1_e0[36] ), 
          .S1(\nZ1_e0[37] ));
    defparam add_952_22.INIT0 = 16'h5666;
    defparam add_952_22.INIT1 = 16'h5666;
    defparam add_952_22.INJECT1_0 = "NO";
    defparam add_952_22.INJECT1_1 = "NO";
    CCU2D add_952_20 (.A0(buf_x[1902]), .B0(buf_x[1931]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1903]), .B1(buf_x[1932]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62147), .COUT(n62148), .S0(\nZ1_e0[34] ), 
          .S1(\nZ1_e0[35] ));
    defparam add_952_20.INIT0 = 16'h5666;
    defparam add_952_20.INIT1 = 16'h5666;
    defparam add_952_20.INJECT1_0 = "NO";
    defparam add_952_20.INJECT1_1 = "NO";
    CCU2D add_952_18 (.A0(buf_x[1900]), .B0(buf_x[1929]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1901]), .B1(buf_x[1930]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62146), .COUT(n62147), .S0(\nZ1_e0[32] ), 
          .S1(\nZ1_e0[33] ));
    defparam add_952_18.INIT0 = 16'h5666;
    defparam add_952_18.INIT1 = 16'h5666;
    defparam add_952_18.INJECT1_0 = "NO";
    defparam add_952_18.INJECT1_1 = "NO";
    CCU2D add_952_16 (.A0(buf_x[1898]), .B0(buf_x[1927]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1899]), .B1(buf_x[1928]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62145), .COUT(n62146), .S0(\nZ1_e0[30] ), 
          .S1(\nZ1_e0[31] ));
    defparam add_952_16.INIT0 = 16'h5666;
    defparam add_952_16.INIT1 = 16'h5666;
    defparam add_952_16.INJECT1_0 = "NO";
    defparam add_952_16.INJECT1_1 = "NO";
    CCU2D add_952_14 (.A0(buf_x[1896]), .B0(buf_x[1925]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1897]), .B1(buf_x[1926]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62144), .COUT(n62145), .S1(\nZ1_e0[29] ));
    defparam add_952_14.INIT0 = 16'h5666;
    defparam add_952_14.INIT1 = 16'h5666;
    defparam add_952_14.INJECT1_0 = "NO";
    defparam add_952_14.INJECT1_1 = "NO";
    CCU2D add_952_12 (.A0(buf_x[1894]), .B0(buf_x[1923]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1895]), .B1(buf_x[1924]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62143), .COUT(n62144));
    defparam add_952_12.INIT0 = 16'h5666;
    defparam add_952_12.INIT1 = 16'h5666;
    defparam add_952_12.INJECT1_0 = "NO";
    defparam add_952_12.INJECT1_1 = "NO";
    CCU2D add_952_10 (.A0(buf_x[1892]), .B0(buf_x[1921]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1893]), .B1(buf_x[1922]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62142), .COUT(n62143));
    defparam add_952_10.INIT0 = 16'h5666;
    defparam add_952_10.INIT1 = 16'h5666;
    defparam add_952_10.INJECT1_0 = "NO";
    defparam add_952_10.INJECT1_1 = "NO";
    CCU2D add_952_8 (.A0(buf_x[1890]), .B0(buf_x[1919]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1891]), .B1(buf_x[1920]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62141), .COUT(n62142));
    defparam add_952_8.INIT0 = 16'h5666;
    defparam add_952_8.INIT1 = 16'h5666;
    defparam add_952_8.INJECT1_0 = "NO";
    defparam add_952_8.INJECT1_1 = "NO";
    CCU2D add_952_6 (.A0(buf_x[1888]), .B0(buf_x[1917]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1889]), .B1(buf_x[1918]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62140), .COUT(n62141));
    defparam add_952_6.INIT0 = 16'h5666;
    defparam add_952_6.INIT1 = 16'h5666;
    defparam add_952_6.INJECT1_0 = "NO";
    defparam add_952_6.INJECT1_1 = "NO";
    CCU2D add_952_4 (.A0(buf_x[1886]), .B0(buf_x[1915]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1887]), .B1(buf_x[1916]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62139), .COUT(n62140));
    defparam add_952_4.INIT0 = 16'h5666;
    defparam add_952_4.INIT1 = 16'h5666;
    defparam add_952_4.INJECT1_0 = "NO";
    defparam add_952_4.INJECT1_1 = "NO";
    CCU2D add_952_2 (.A0(buf_x[1884]), .B0(buf_x[1913]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1885]), .B1(buf_x[1914]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62139));
    defparam add_952_2.INIT0 = 16'h7000;
    defparam add_952_2.INIT1 = 16'h5666;
    defparam add_952_2.INJECT1_0 = "NO";
    defparam add_952_2.INJECT1_1 = "NO";
    CCU2D add_496_38 (.A0(buf_r[1756]), .B0(buf_r[1793]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62138), .S0(buf_x[1912]));
    defparam add_496_38.INIT0 = 16'h5666;
    defparam add_496_38.INIT1 = 16'h0000;
    defparam add_496_38.INJECT1_0 = "NO";
    defparam add_496_38.INJECT1_1 = "NO";
    CCU2D add_496_36 (.A0(buf_r[1756]), .B0(buf_r[1791]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1756]), .B1(buf_r[1792]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62137), .COUT(n62138), .S0(buf_x[1910]), 
          .S1(buf_x[1911]));
    defparam add_496_36.INIT0 = 16'h5666;
    defparam add_496_36.INIT1 = 16'h5666;
    defparam add_496_36.INJECT1_0 = "NO";
    defparam add_496_36.INJECT1_1 = "NO";
    CCU2D add_496_34 (.A0(buf_r[1756]), .B0(buf_r[1789]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1756]), .B1(buf_r[1790]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62136), .COUT(n62137), .S0(buf_x[1908]), 
          .S1(buf_x[1909]));
    defparam add_496_34.INIT0 = 16'h5666;
    defparam add_496_34.INIT1 = 16'h5666;
    defparam add_496_34.INJECT1_0 = "NO";
    defparam add_496_34.INJECT1_1 = "NO";
    CCU2D add_496_32 (.A0(buf_r[1756]), .B0(buf_r[1787]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1756]), .B1(buf_r[1788]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62135), .COUT(n62136), .S0(buf_x[1906]), 
          .S1(buf_x[1907]));
    defparam add_496_32.INIT0 = 16'h5666;
    defparam add_496_32.INIT1 = 16'h5666;
    defparam add_496_32.INJECT1_0 = "NO";
    defparam add_496_32.INJECT1_1 = "NO";
    CCU2D add_496_30 (.A0(buf_r[1756]), .B0(buf_r[1785]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1756]), .B1(buf_r[1786]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62134), .COUT(n62135), .S0(buf_x[1904]), 
          .S1(buf_x[1905]));
    defparam add_496_30.INIT0 = 16'h5666;
    defparam add_496_30.INIT1 = 16'h5666;
    defparam add_496_30.INJECT1_0 = "NO";
    defparam add_496_30.INJECT1_1 = "NO";
    CCU2D add_496_28 (.A0(buf_r[1754]), .B0(buf_r[1783]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1755]), .B1(buf_r[1784]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62133), .COUT(n62134), .S0(buf_x[1902]), 
          .S1(buf_x[1903]));
    defparam add_496_28.INIT0 = 16'h5666;
    defparam add_496_28.INIT1 = 16'h5666;
    defparam add_496_28.INJECT1_0 = "NO";
    defparam add_496_28.INJECT1_1 = "NO";
    CCU2D add_496_26 (.A0(buf_r[1752]), .B0(buf_r[1781]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1753]), .B1(buf_r[1782]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62132), .COUT(n62133), .S0(buf_x[1900]), 
          .S1(buf_x[1901]));
    defparam add_496_26.INIT0 = 16'h5666;
    defparam add_496_26.INIT1 = 16'h5666;
    defparam add_496_26.INJECT1_0 = "NO";
    defparam add_496_26.INJECT1_1 = "NO";
    CCU2D add_496_24 (.A0(buf_r[1750]), .B0(buf_r[1779]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1751]), .B1(buf_r[1780]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62131), .COUT(n62132), .S0(buf_x[1898]), 
          .S1(buf_x[1899]));
    defparam add_496_24.INIT0 = 16'h5666;
    defparam add_496_24.INIT1 = 16'h5666;
    defparam add_496_24.INJECT1_0 = "NO";
    defparam add_496_24.INJECT1_1 = "NO";
    CCU2D add_496_22 (.A0(buf_r[1748]), .B0(buf_r[1777]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1749]), .B1(buf_r[1778]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62130), .COUT(n62131), .S0(buf_x[1896]), 
          .S1(buf_x[1897]));
    defparam add_496_22.INIT0 = 16'h5666;
    defparam add_496_22.INIT1 = 16'h5666;
    defparam add_496_22.INJECT1_0 = "NO";
    defparam add_496_22.INJECT1_1 = "NO";
    CCU2D add_496_20 (.A0(buf_r[1746]), .B0(buf_r[1775]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1747]), .B1(buf_r[1776]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62129), .COUT(n62130), .S0(buf_x[1894]), 
          .S1(buf_x[1895]));
    defparam add_496_20.INIT0 = 16'h5666;
    defparam add_496_20.INIT1 = 16'h5666;
    defparam add_496_20.INJECT1_0 = "NO";
    defparam add_496_20.INJECT1_1 = "NO";
    CCU2D add_496_18 (.A0(buf_r[1744]), .B0(buf_r[1773]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1745]), .B1(buf_r[1774]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62128), .COUT(n62129), .S0(buf_x[1892]), 
          .S1(buf_x[1893]));
    defparam add_496_18.INIT0 = 16'h5666;
    defparam add_496_18.INIT1 = 16'h5666;
    defparam add_496_18.INJECT1_0 = "NO";
    defparam add_496_18.INJECT1_1 = "NO";
    CCU2D add_496_16 (.A0(buf_r[1742]), .B0(buf_r[1771]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1743]), .B1(buf_r[1772]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62127), .COUT(n62128), .S0(buf_x[1890]), 
          .S1(buf_x[1891]));
    defparam add_496_16.INIT0 = 16'h5666;
    defparam add_496_16.INIT1 = 16'h5666;
    defparam add_496_16.INJECT1_0 = "NO";
    defparam add_496_16.INJECT1_1 = "NO";
    CCU2D add_496_14 (.A0(buf_r[1740]), .B0(buf_r[1769]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1741]), .B1(buf_r[1770]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62126), .COUT(n62127), .S0(buf_x[1888]), 
          .S1(buf_x[1889]));
    defparam add_496_14.INIT0 = 16'h5666;
    defparam add_496_14.INIT1 = 16'h5666;
    defparam add_496_14.INJECT1_0 = "NO";
    defparam add_496_14.INJECT1_1 = "NO";
    CCU2D add_496_12 (.A0(buf_r[1738]), .B0(buf_r[1767]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1739]), .B1(buf_r[1768]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62125), .COUT(n62126), .S0(buf_x[1886]), 
          .S1(buf_x[1887]));
    defparam add_496_12.INIT0 = 16'h5666;
    defparam add_496_12.INIT1 = 16'h5666;
    defparam add_496_12.INJECT1_0 = "NO";
    defparam add_496_12.INJECT1_1 = "NO";
    CCU2D add_496_10 (.A0(buf_r[1736]), .B0(buf_r[1765]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1737]), .B1(buf_r[1766]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62124), .COUT(n62125), .S0(buf_x[1884]), 
          .S1(buf_x[1885]));
    defparam add_496_10.INIT0 = 16'h5666;
    defparam add_496_10.INIT1 = 16'h5666;
    defparam add_496_10.INJECT1_0 = "NO";
    defparam add_496_10.INJECT1_1 = "NO";
    CCU2D add_496_8 (.A0(buf_r[1734]), .B0(buf_r[1763]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1735]), .B1(buf_r[1764]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62123), .COUT(n62124));
    defparam add_496_8.INIT0 = 16'h5666;
    defparam add_496_8.INIT1 = 16'h5666;
    defparam add_496_8.INJECT1_0 = "NO";
    defparam add_496_8.INJECT1_1 = "NO";
    CCU2D add_496_6 (.A0(buf_r[1732]), .B0(buf_r[1761]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1733]), .B1(buf_r[1762]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62122), .COUT(n62123));
    defparam add_496_6.INIT0 = 16'h5666;
    defparam add_496_6.INIT1 = 16'h5666;
    defparam add_496_6.INJECT1_0 = "NO";
    defparam add_496_6.INJECT1_1 = "NO";
    CCU2D add_496_4 (.A0(buf_r[1730]), .B0(buf_r[1759]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1731]), .B1(buf_r[1760]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62121), .COUT(n62122));
    defparam add_496_4.INIT0 = 16'h5666;
    defparam add_496_4.INIT1 = 16'h5666;
    defparam add_496_4.INJECT1_0 = "NO";
    defparam add_496_4.INJECT1_1 = "NO";
    CCU2D add_496_2 (.A0(buf_r[1728]), .B0(buf_r[1757]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1729]), .B1(buf_r[1758]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62121));
    defparam add_496_2.INIT0 = 16'h7000;
    defparam add_496_2.INIT1 = 16'h5666;
    defparam add_496_2.INJECT1_0 = "NO";
    defparam add_496_2.INJECT1_1 = "NO";
    CCU2D add_383_34 (.A0(buf_x[1554]), .B0(buf_x[1587]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62116), .S0(buf_x[1793]));
    defparam add_383_34.INIT0 = 16'h5666;
    defparam add_383_34.INIT1 = 16'h0000;
    defparam add_383_34.INJECT1_0 = "NO";
    defparam add_383_34.INJECT1_1 = "NO";
    CCU2D add_383_32 (.A0(buf_x[1554]), .B0(buf_x[1585]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1554]), .B1(buf_x[1586]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62115), .COUT(n62116), .S0(buf_x[1791]), 
          .S1(buf_x[1792]));
    defparam add_383_32.INIT0 = 16'h5666;
    defparam add_383_32.INIT1 = 16'h5666;
    defparam add_383_32.INJECT1_0 = "NO";
    defparam add_383_32.INJECT1_1 = "NO";
    CCU2D add_383_30 (.A0(buf_x[1554]), .B0(buf_x[1583]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1554]), .B1(buf_x[1584]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62114), .COUT(n62115), .S0(buf_x[1789]), 
          .S1(buf_x[1790]));
    defparam add_383_30.INIT0 = 16'h5666;
    defparam add_383_30.INIT1 = 16'h5666;
    defparam add_383_30.INJECT1_0 = "NO";
    defparam add_383_30.INJECT1_1 = "NO";
    CCU2D add_383_28 (.A0(buf_x[1552]), .B0(buf_x[1581]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1553]), .B1(buf_x[1582]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62113), .COUT(n62114), .S0(buf_x[1787]), 
          .S1(buf_x[1788]));
    defparam add_383_28.INIT0 = 16'h5666;
    defparam add_383_28.INIT1 = 16'h5666;
    defparam add_383_28.INJECT1_0 = "NO";
    defparam add_383_28.INJECT1_1 = "NO";
    CCU2D add_383_26 (.A0(buf_x[1550]), .B0(buf_x[1579]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1551]), .B1(buf_x[1580]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62112), .COUT(n62113), .S0(buf_x[1785]), 
          .S1(buf_x[1786]));
    defparam add_383_26.INIT0 = 16'h5666;
    defparam add_383_26.INIT1 = 16'h5666;
    defparam add_383_26.INJECT1_0 = "NO";
    defparam add_383_26.INJECT1_1 = "NO";
    CCU2D add_383_24 (.A0(buf_x[1548]), .B0(buf_x[1577]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1549]), .B1(buf_x[1578]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62111), .COUT(n62112), .S0(buf_x[1783]), 
          .S1(buf_x[1784]));
    defparam add_383_24.INIT0 = 16'h5666;
    defparam add_383_24.INIT1 = 16'h5666;
    defparam add_383_24.INJECT1_0 = "NO";
    defparam add_383_24.INJECT1_1 = "NO";
    CCU2D add_383_22 (.A0(buf_x[1546]), .B0(buf_x[1575]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1547]), .B1(buf_x[1576]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62110), .COUT(n62111), .S0(buf_x[1781]), 
          .S1(buf_x[1782]));
    defparam add_383_22.INIT0 = 16'h5666;
    defparam add_383_22.INIT1 = 16'h5666;
    defparam add_383_22.INJECT1_0 = "NO";
    defparam add_383_22.INJECT1_1 = "NO";
    CCU2D add_383_20 (.A0(buf_x[1544]), .B0(buf_x[1573]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1545]), .B1(buf_x[1574]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62109), .COUT(n62110), .S0(buf_x[1779]), 
          .S1(buf_x[1780]));
    defparam add_383_20.INIT0 = 16'h5666;
    defparam add_383_20.INIT1 = 16'h5666;
    defparam add_383_20.INJECT1_0 = "NO";
    defparam add_383_20.INJECT1_1 = "NO";
    CCU2D add_383_18 (.A0(buf_x[1542]), .B0(buf_x[1571]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1543]), .B1(buf_x[1572]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62108), .COUT(n62109), .S0(buf_x[1777]), 
          .S1(buf_x[1778]));
    defparam add_383_18.INIT0 = 16'h5666;
    defparam add_383_18.INIT1 = 16'h5666;
    defparam add_383_18.INJECT1_0 = "NO";
    defparam add_383_18.INJECT1_1 = "NO";
    CCU2D add_383_16 (.A0(buf_x[1540]), .B0(buf_x[1569]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1541]), .B1(buf_x[1570]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62107), .COUT(n62108), .S0(buf_x[1775]), 
          .S1(buf_x[1776]));
    defparam add_383_16.INIT0 = 16'h5666;
    defparam add_383_16.INIT1 = 16'h5666;
    defparam add_383_16.INJECT1_0 = "NO";
    defparam add_383_16.INJECT1_1 = "NO";
    CCU2D add_383_14 (.A0(buf_x[1538]), .B0(buf_x[1567]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1539]), .B1(buf_x[1568]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62106), .COUT(n62107), .S0(buf_x[1773]), 
          .S1(buf_x[1774]));
    defparam add_383_14.INIT0 = 16'h5666;
    defparam add_383_14.INIT1 = 16'h5666;
    defparam add_383_14.INJECT1_0 = "NO";
    defparam add_383_14.INJECT1_1 = "NO";
    CCU2D add_383_12 (.A0(buf_x[1536]), .B0(buf_x[1565]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1537]), .B1(buf_x[1566]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62105), .COUT(n62106), .S0(buf_x[1771]), 
          .S1(buf_x[1772]));
    defparam add_383_12.INIT0 = 16'h5666;
    defparam add_383_12.INIT1 = 16'h5666;
    defparam add_383_12.INJECT1_0 = "NO";
    defparam add_383_12.INJECT1_1 = "NO";
    CCU2D add_383_10 (.A0(buf_x[1534]), .B0(buf_x[1563]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1535]), .B1(buf_x[1564]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62104), .COUT(n62105), .S0(buf_x[1769]), 
          .S1(buf_x[1770]));
    defparam add_383_10.INIT0 = 16'h5666;
    defparam add_383_10.INIT1 = 16'h5666;
    defparam add_383_10.INJECT1_0 = "NO";
    defparam add_383_10.INJECT1_1 = "NO";
    CCU2D add_383_8 (.A0(buf_x[1532]), .B0(buf_x[1561]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1533]), .B1(buf_x[1562]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62103), .COUT(n62104), .S0(buf_x[1767]), 
          .S1(buf_x[1768]));
    defparam add_383_8.INIT0 = 16'h5666;
    defparam add_383_8.INIT1 = 16'h5666;
    defparam add_383_8.INJECT1_0 = "NO";
    defparam add_383_8.INJECT1_1 = "NO";
    CCU2D add_383_6 (.A0(buf_x[1530]), .B0(buf_x[1559]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1531]), .B1(buf_x[1560]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62102), .COUT(n62103), .S0(buf_x[1765]), 
          .S1(buf_x[1766]));
    defparam add_383_6.INIT0 = 16'h5666;
    defparam add_383_6.INIT1 = 16'h5666;
    defparam add_383_6.INJECT1_0 = "NO";
    defparam add_383_6.INJECT1_1 = "NO";
    CCU2D add_383_4 (.A0(buf_r[1148]), .B0(buf_r[1177]), .C0(buf_x[1528]), 
          .D0(GND_net), .A1(buf_x[1529]), .B1(buf_x[1558]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62101), .COUT(n62102), .S0(buf_x[1763]), 
          .S1(buf_x[1764]));
    defparam add_383_4.INIT0 = 16'h9696;
    defparam add_383_4.INIT1 = 16'h5666;
    defparam add_383_4.INJECT1_0 = "NO";
    defparam add_383_4.INJECT1_1 = "NO";
    CCU2D add_383_2 (.A0(buf_x[1526]), .B0(buf_x[1555]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1527]), .B1(buf_x[1556]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62101), .S1(buf_x[1762]));
    defparam add_383_2.INIT0 = 16'h7000;
    defparam add_383_2.INIT1 = 16'h5666;
    defparam add_383_2.INJECT1_0 = "NO";
    defparam add_383_2.INJECT1_1 = "NO";
    CCU2D add_382_34 (.A0(buf_x[1488]), .B0(buf_x[1521]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62099), .S0(buf_x[1756]));
    defparam add_382_34.INIT0 = 16'h5666;
    defparam add_382_34.INIT1 = 16'h0000;
    defparam add_382_34.INJECT1_0 = "NO";
    defparam add_382_34.INJECT1_1 = "NO";
    CCU2D add_382_32 (.A0(buf_x[1488]), .B0(buf_x[1519]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1488]), .B1(buf_x[1520]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62098), .COUT(n62099), .S0(buf_x[1754]), 
          .S1(buf_x[1755]));
    defparam add_382_32.INIT0 = 16'h5666;
    defparam add_382_32.INIT1 = 16'h5666;
    defparam add_382_32.INJECT1_0 = "NO";
    defparam add_382_32.INJECT1_1 = "NO";
    CCU2D add_382_30 (.A0(buf_x[1488]), .B0(buf_x[1517]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1488]), .B1(buf_x[1518]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62097), .COUT(n62098), .S0(buf_x[1752]), 
          .S1(buf_x[1753]));
    defparam add_382_30.INIT0 = 16'h5666;
    defparam add_382_30.INIT1 = 16'h5666;
    defparam add_382_30.INJECT1_0 = "NO";
    defparam add_382_30.INJECT1_1 = "NO";
    CCU2D add_382_28 (.A0(buf_x[1486]), .B0(buf_x[1515]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1487]), .B1(buf_x[1516]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62096), .COUT(n62097), .S0(buf_x[1750]), 
          .S1(buf_x[1751]));
    defparam add_382_28.INIT0 = 16'h5666;
    defparam add_382_28.INIT1 = 16'h5666;
    defparam add_382_28.INJECT1_0 = "NO";
    defparam add_382_28.INJECT1_1 = "NO";
    CCU2D add_382_26 (.A0(buf_x[1484]), .B0(buf_x[1513]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1485]), .B1(buf_x[1514]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62095), .COUT(n62096), .S0(buf_x[1748]), 
          .S1(buf_x[1749]));
    defparam add_382_26.INIT0 = 16'h5666;
    defparam add_382_26.INIT1 = 16'h5666;
    defparam add_382_26.INJECT1_0 = "NO";
    defparam add_382_26.INJECT1_1 = "NO";
    CCU2D add_382_24 (.A0(buf_x[1482]), .B0(buf_x[1511]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1483]), .B1(buf_x[1512]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62094), .COUT(n62095), .S0(buf_x[1746]), 
          .S1(buf_x[1747]));
    defparam add_382_24.INIT0 = 16'h5666;
    defparam add_382_24.INIT1 = 16'h5666;
    defparam add_382_24.INJECT1_0 = "NO";
    defparam add_382_24.INJECT1_1 = "NO";
    CCU2D add_382_22 (.A0(buf_x[1480]), .B0(buf_x[1509]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1481]), .B1(buf_x[1510]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62093), .COUT(n62094), .S0(buf_x[1744]), 
          .S1(buf_x[1745]));
    defparam add_382_22.INIT0 = 16'h5666;
    defparam add_382_22.INIT1 = 16'h5666;
    defparam add_382_22.INJECT1_0 = "NO";
    defparam add_382_22.INJECT1_1 = "NO";
    CCU2D add_382_20 (.A0(buf_x[1478]), .B0(buf_x[1507]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1479]), .B1(buf_x[1508]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62092), .COUT(n62093), .S0(buf_x[1742]), 
          .S1(buf_x[1743]));
    defparam add_382_20.INIT0 = 16'h5666;
    defparam add_382_20.INIT1 = 16'h5666;
    defparam add_382_20.INJECT1_0 = "NO";
    defparam add_382_20.INJECT1_1 = "NO";
    CCU2D add_382_18 (.A0(buf_x[1476]), .B0(buf_x[1505]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1477]), .B1(buf_x[1506]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62091), .COUT(n62092), .S0(buf_x[1740]), 
          .S1(buf_x[1741]));
    defparam add_382_18.INIT0 = 16'h5666;
    defparam add_382_18.INIT1 = 16'h5666;
    defparam add_382_18.INJECT1_0 = "NO";
    defparam add_382_18.INJECT1_1 = "NO";
    CCU2D add_382_16 (.A0(buf_x[1474]), .B0(buf_x[1503]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1475]), .B1(buf_x[1504]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62090), .COUT(n62091), .S0(buf_x[1738]), 
          .S1(buf_x[1739]));
    defparam add_382_16.INIT0 = 16'h5666;
    defparam add_382_16.INIT1 = 16'h5666;
    defparam add_382_16.INJECT1_0 = "NO";
    defparam add_382_16.INJECT1_1 = "NO";
    CCU2D add_382_14 (.A0(buf_x[1472]), .B0(buf_x[1501]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1473]), .B1(buf_x[1502]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62089), .COUT(n62090), .S0(buf_x[1736]), 
          .S1(buf_x[1737]));
    defparam add_382_14.INIT0 = 16'h5666;
    defparam add_382_14.INIT1 = 16'h5666;
    defparam add_382_14.INJECT1_0 = "NO";
    defparam add_382_14.INJECT1_1 = "NO";
    CCU2D add_382_12 (.A0(buf_x[1470]), .B0(buf_x[1499]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1471]), .B1(buf_x[1500]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62088), .COUT(n62089), .S0(buf_x[1734]), 
          .S1(buf_x[1735]));
    defparam add_382_12.INIT0 = 16'h5666;
    defparam add_382_12.INIT1 = 16'h5666;
    defparam add_382_12.INJECT1_0 = "NO";
    defparam add_382_12.INJECT1_1 = "NO";
    CCU2D add_382_10 (.A0(buf_x[1468]), .B0(buf_x[1497]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1469]), .B1(buf_x[1498]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62087), .COUT(n62088), .S0(buf_x[1732]), 
          .S1(buf_x[1733]));
    defparam add_382_10.INIT0 = 16'h5666;
    defparam add_382_10.INIT1 = 16'h5666;
    defparam add_382_10.INJECT1_0 = "NO";
    defparam add_382_10.INJECT1_1 = "NO";
    CCU2D add_382_8 (.A0(buf_x[1466]), .B0(buf_x[1495]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1467]), .B1(buf_x[1496]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62086), .COUT(n62087), .S0(buf_x[1730]), 
          .S1(buf_x[1731]));
    defparam add_382_8.INIT0 = 16'h5666;
    defparam add_382_8.INIT1 = 16'h5666;
    defparam add_382_8.INJECT1_0 = "NO";
    defparam add_382_8.INJECT1_1 = "NO";
    CCU2D add_382_6 (.A0(buf_x[1464]), .B0(buf_x[1493]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1465]), .B1(buf_x[1494]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62085), .COUT(n62086), .S0(buf_x[1728]), 
          .S1(buf_x[1729]));
    defparam add_382_6.INIT0 = 16'h5666;
    defparam add_382_6.INIT1 = 16'h5666;
    defparam add_382_6.INJECT1_0 = "NO";
    defparam add_382_6.INJECT1_1 = "NO";
    CCU2D add_382_4 (.A0(buf_r[1024]), .B0(buf_r[1053]), .C0(buf_x[1462]), 
          .D0(GND_net), .A1(buf_x[1463]), .B1(buf_x[1492]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62084), .COUT(n62085));
    defparam add_382_4.INIT0 = 16'h9696;
    defparam add_382_4.INIT1 = 16'h5666;
    defparam add_382_4.INJECT1_0 = "NO";
    defparam add_382_4.INJECT1_1 = "NO";
    CCU2D add_382_2 (.A0(buf_x[1460]), .B0(buf_x[1489]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1461]), .B1(buf_x[1490]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62084));
    defparam add_382_2.INIT0 = 16'h7000;
    defparam add_382_2.INIT1 = 16'h5666;
    defparam add_382_2.INJECT1_0 = "NO";
    defparam add_382_2.INJECT1_1 = "NO";
    CCU2D add_4618_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62079), 
          .S0(buf_x[1620]));
    defparam add_4618_cout.INIT0 = 16'h0000;
    defparam add_4618_cout.INIT1 = 16'h0000;
    defparam add_4618_cout.INJECT1_0 = "NO";
    defparam add_4618_cout.INJECT1_1 = "NO";
    CCU2D add_4618_30 (.A0(buf_r[1267]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_r[1268]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62078), .COUT(n62079), .S0(buf_x[1618]), .S1(buf_x[1619]));
    defparam add_4618_30.INIT0 = 16'hfaaa;
    defparam add_4618_30.INIT1 = 16'hfaaa;
    defparam add_4618_30.INJECT1_0 = "NO";
    defparam add_4618_30.INJECT1_1 = "NO";
    CCU2D add_4618_28 (.A0(buf_r[1236]), .B0(buf_r[1265]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1237]), .B1(buf_r[1266]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62077), .COUT(n62078), .S0(buf_x[1616]), 
          .S1(buf_x[1617]));
    defparam add_4618_28.INIT0 = 16'h5666;
    defparam add_4618_28.INIT1 = 16'h5666;
    defparam add_4618_28.INJECT1_0 = "NO";
    defparam add_4618_28.INJECT1_1 = "NO";
    CCU2D add_4618_26 (.A0(buf_r[1234]), .B0(buf_r[1263]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1235]), .B1(buf_r[1264]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62076), .COUT(n62077), .S0(buf_x[1614]), 
          .S1(buf_x[1615]));
    defparam add_4618_26.INIT0 = 16'h5666;
    defparam add_4618_26.INIT1 = 16'h5666;
    defparam add_4618_26.INJECT1_0 = "NO";
    defparam add_4618_26.INJECT1_1 = "NO";
    CCU2D add_4618_24 (.A0(buf_r[1232]), .B0(buf_r[1261]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1233]), .B1(buf_r[1262]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62075), .COUT(n62076), .S0(buf_x[1612]), 
          .S1(buf_x[1613]));
    defparam add_4618_24.INIT0 = 16'h5666;
    defparam add_4618_24.INIT1 = 16'h5666;
    defparam add_4618_24.INJECT1_0 = "NO";
    defparam add_4618_24.INJECT1_1 = "NO";
    CCU2D add_4618_22 (.A0(buf_r[1230]), .B0(buf_r[1259]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1231]), .B1(buf_r[1260]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62074), .COUT(n62075), .S0(buf_x[1610]), 
          .S1(buf_x[1611]));
    defparam add_4618_22.INIT0 = 16'h5666;
    defparam add_4618_22.INIT1 = 16'h5666;
    defparam add_4618_22.INJECT1_0 = "NO";
    defparam add_4618_22.INJECT1_1 = "NO";
    CCU2D add_4618_20 (.A0(buf_r[1228]), .B0(buf_r[1257]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1229]), .B1(buf_r[1258]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62073), .COUT(n62074), .S0(buf_x[1608]), 
          .S1(buf_x[1609]));
    defparam add_4618_20.INIT0 = 16'h5666;
    defparam add_4618_20.INIT1 = 16'h5666;
    defparam add_4618_20.INJECT1_0 = "NO";
    defparam add_4618_20.INJECT1_1 = "NO";
    CCU2D add_4618_18 (.A0(buf_r[1226]), .B0(buf_r[1255]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1227]), .B1(buf_r[1256]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62072), .COUT(n62073), .S0(buf_x[1606]), 
          .S1(buf_x[1607]));
    defparam add_4618_18.INIT0 = 16'h5666;
    defparam add_4618_18.INIT1 = 16'h5666;
    defparam add_4618_18.INJECT1_0 = "NO";
    defparam add_4618_18.INJECT1_1 = "NO";
    CCU2D add_4618_16 (.A0(buf_r[1224]), .B0(buf_r[1253]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1225]), .B1(buf_r[1254]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62071), .COUT(n62072), .S0(buf_x[1604]), 
          .S1(buf_x[1605]));
    defparam add_4618_16.INIT0 = 16'h5666;
    defparam add_4618_16.INIT1 = 16'h5666;
    defparam add_4618_16.INJECT1_0 = "NO";
    defparam add_4618_16.INJECT1_1 = "NO";
    CCU2D add_4618_14 (.A0(buf_r[1222]), .B0(buf_r[1251]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1223]), .B1(buf_r[1252]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62070), .COUT(n62071), .S0(buf_x[1602]), 
          .S1(buf_x[1603]));
    defparam add_4618_14.INIT0 = 16'h5666;
    defparam add_4618_14.INIT1 = 16'h5666;
    defparam add_4618_14.INJECT1_0 = "NO";
    defparam add_4618_14.INJECT1_1 = "NO";
    CCU2D add_4618_12 (.A0(buf_r[1220]), .B0(buf_r[1249]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1221]), .B1(buf_r[1250]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62069), .COUT(n62070), .S0(buf_x[1600]), 
          .S1(buf_x[1601]));
    defparam add_4618_12.INIT0 = 16'h5666;
    defparam add_4618_12.INIT1 = 16'h5666;
    defparam add_4618_12.INJECT1_0 = "NO";
    defparam add_4618_12.INJECT1_1 = "NO";
    CCU2D add_4618_10 (.A0(buf_r[1218]), .B0(buf_r[1247]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1219]), .B1(buf_r[1248]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62068), .COUT(n62069), .S0(buf_x[1598]), 
          .S1(buf_x[1599]));
    defparam add_4618_10.INIT0 = 16'h5666;
    defparam add_4618_10.INIT1 = 16'h5666;
    defparam add_4618_10.INJECT1_0 = "NO";
    defparam add_4618_10.INJECT1_1 = "NO";
    CCU2D add_4618_8 (.A0(buf_r[1216]), .B0(buf_r[1245]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1217]), .B1(buf_r[1246]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62067), .COUT(n62068), .S0(buf_x[1596]), 
          .S1(buf_x[1597]));
    defparam add_4618_8.INIT0 = 16'h5666;
    defparam add_4618_8.INIT1 = 16'h5666;
    defparam add_4618_8.INJECT1_0 = "NO";
    defparam add_4618_8.INJECT1_1 = "NO";
    CCU2D add_4618_6 (.A0(buf_r[1214]), .B0(buf_r[1243]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1215]), .B1(buf_r[1244]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62066), .COUT(n62067), .S0(buf_x[1594]), 
          .S1(buf_x[1595]));
    defparam add_4618_6.INIT0 = 16'h5666;
    defparam add_4618_6.INIT1 = 16'h5666;
    defparam add_4618_6.INJECT1_0 = "NO";
    defparam add_4618_6.INJECT1_1 = "NO";
    CCU2D add_4618_4 (.A0(buf_r[1212]), .B0(buf_r[1241]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1213]), .B1(buf_r[1242]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62065), .COUT(n62066), .S0(buf_x[1592]), 
          .S1(buf_x[1593]));
    defparam add_4618_4.INIT0 = 16'h5666;
    defparam add_4618_4.INIT1 = 16'h5666;
    defparam add_4618_4.INJECT1_0 = "NO";
    defparam add_4618_4.INJECT1_1 = "NO";
    CCU2D add_4618_2 (.A0(buf_r[1210]), .B0(buf_r[1239]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1211]), .B1(buf_r[1240]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62065), .S1(buf_x[1797]));
    defparam add_4618_2.INIT0 = 16'h7000;
    defparam add_4618_2.INIT1 = 16'h5666;
    defparam add_4618_2.INJECT1_0 = "NO";
    defparam add_4618_2.INJECT1_1 = "NO";
    CCU2D add_4617_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62063), 
          .S0(buf_x[1587]));
    defparam add_4617_cout.INIT0 = 16'h0000;
    defparam add_4617_cout.INIT1 = 16'h0000;
    defparam add_4617_cout.INJECT1_0 = "NO";
    defparam add_4617_cout.INJECT1_1 = "NO";
    CCU2D add_4617_30 (.A0(buf_r[1205]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_r[1206]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62062), .COUT(n62063), .S0(buf_x[1585]), .S1(buf_x[1586]));
    defparam add_4617_30.INIT0 = 16'hfaaa;
    defparam add_4617_30.INIT1 = 16'hfaaa;
    defparam add_4617_30.INJECT1_0 = "NO";
    defparam add_4617_30.INJECT1_1 = "NO";
    CCU2D add_4617_28 (.A0(buf_r[1174]), .B0(buf_r[1203]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1175]), .B1(buf_r[1204]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62061), .COUT(n62062), .S0(buf_x[1583]), 
          .S1(buf_x[1584]));
    defparam add_4617_28.INIT0 = 16'h5666;
    defparam add_4617_28.INIT1 = 16'h5666;
    defparam add_4617_28.INJECT1_0 = "NO";
    defparam add_4617_28.INJECT1_1 = "NO";
    CCU2D add_4617_26 (.A0(buf_r[1172]), .B0(buf_r[1201]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1173]), .B1(buf_r[1202]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62060), .COUT(n62061), .S0(buf_x[1581]), 
          .S1(buf_x[1582]));
    defparam add_4617_26.INIT0 = 16'h5666;
    defparam add_4617_26.INIT1 = 16'h5666;
    defparam add_4617_26.INJECT1_0 = "NO";
    defparam add_4617_26.INJECT1_1 = "NO";
    CCU2D add_4617_24 (.A0(buf_r[1170]), .B0(buf_r[1199]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1171]), .B1(buf_r[1200]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62059), .COUT(n62060), .S0(buf_x[1579]), 
          .S1(buf_x[1580]));
    defparam add_4617_24.INIT0 = 16'h5666;
    defparam add_4617_24.INIT1 = 16'h5666;
    defparam add_4617_24.INJECT1_0 = "NO";
    defparam add_4617_24.INJECT1_1 = "NO";
    CCU2D add_4617_22 (.A0(buf_r[1168]), .B0(buf_r[1197]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1169]), .B1(buf_r[1198]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62058), .COUT(n62059), .S0(buf_x[1577]), 
          .S1(buf_x[1578]));
    defparam add_4617_22.INIT0 = 16'h5666;
    defparam add_4617_22.INIT1 = 16'h5666;
    defparam add_4617_22.INJECT1_0 = "NO";
    defparam add_4617_22.INJECT1_1 = "NO";
    CCU2D add_4617_20 (.A0(buf_r[1166]), .B0(buf_r[1195]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1167]), .B1(buf_r[1196]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62057), .COUT(n62058), .S0(buf_x[1575]), 
          .S1(buf_x[1576]));
    defparam add_4617_20.INIT0 = 16'h5666;
    defparam add_4617_20.INIT1 = 16'h5666;
    defparam add_4617_20.INJECT1_0 = "NO";
    defparam add_4617_20.INJECT1_1 = "NO";
    CCU2D add_4617_18 (.A0(buf_r[1164]), .B0(buf_r[1193]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1165]), .B1(buf_r[1194]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62056), .COUT(n62057), .S0(buf_x[1573]), 
          .S1(buf_x[1574]));
    defparam add_4617_18.INIT0 = 16'h5666;
    defparam add_4617_18.INIT1 = 16'h5666;
    defparam add_4617_18.INJECT1_0 = "NO";
    defparam add_4617_18.INJECT1_1 = "NO";
    CCU2D add_4617_16 (.A0(buf_r[1162]), .B0(buf_r[1191]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1163]), .B1(buf_r[1192]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62055), .COUT(n62056), .S0(buf_x[1571]), 
          .S1(buf_x[1572]));
    defparam add_4617_16.INIT0 = 16'h5666;
    defparam add_4617_16.INIT1 = 16'h5666;
    defparam add_4617_16.INJECT1_0 = "NO";
    defparam add_4617_16.INJECT1_1 = "NO";
    CCU2D add_4617_14 (.A0(buf_r[1160]), .B0(buf_r[1189]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1161]), .B1(buf_r[1190]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62054), .COUT(n62055), .S0(buf_x[1569]), 
          .S1(buf_x[1570]));
    defparam add_4617_14.INIT0 = 16'h5666;
    defparam add_4617_14.INIT1 = 16'h5666;
    defparam add_4617_14.INJECT1_0 = "NO";
    defparam add_4617_14.INJECT1_1 = "NO";
    CCU2D add_4617_12 (.A0(buf_r[1158]), .B0(buf_r[1187]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1159]), .B1(buf_r[1188]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62053), .COUT(n62054), .S0(buf_x[1567]), 
          .S1(buf_x[1568]));
    defparam add_4617_12.INIT0 = 16'h5666;
    defparam add_4617_12.INIT1 = 16'h5666;
    defparam add_4617_12.INJECT1_0 = "NO";
    defparam add_4617_12.INJECT1_1 = "NO";
    CCU2D add_4617_10 (.A0(buf_r[1156]), .B0(buf_r[1185]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1157]), .B1(buf_r[1186]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62052), .COUT(n62053), .S0(buf_x[1565]), 
          .S1(buf_x[1566]));
    defparam add_4617_10.INIT0 = 16'h5666;
    defparam add_4617_10.INIT1 = 16'h5666;
    defparam add_4617_10.INJECT1_0 = "NO";
    defparam add_4617_10.INJECT1_1 = "NO";
    CCU2D add_4617_8 (.A0(buf_r[1154]), .B0(buf_r[1183]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1155]), .B1(buf_r[1184]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62051), .COUT(n62052), .S0(buf_x[1563]), 
          .S1(buf_x[1564]));
    defparam add_4617_8.INIT0 = 16'h5666;
    defparam add_4617_8.INIT1 = 16'h5666;
    defparam add_4617_8.INJECT1_0 = "NO";
    defparam add_4617_8.INJECT1_1 = "NO";
    CCU2D add_4617_6 (.A0(buf_r[1152]), .B0(buf_r[1181]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1153]), .B1(buf_r[1182]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62050), .COUT(n62051), .S0(buf_x[1561]), 
          .S1(buf_x[1562]));
    defparam add_4617_6.INIT0 = 16'h5666;
    defparam add_4617_6.INIT1 = 16'h5666;
    defparam add_4617_6.INJECT1_0 = "NO";
    defparam add_4617_6.INJECT1_1 = "NO";
    CCU2D add_4617_4 (.A0(buf_r[1150]), .B0(buf_r[1179]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1151]), .B1(buf_r[1180]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62049), .COUT(n62050), .S0(buf_x[1559]), 
          .S1(buf_x[1560]));
    defparam add_4617_4.INIT0 = 16'h5666;
    defparam add_4617_4.INIT1 = 16'h5666;
    defparam add_4617_4.INJECT1_0 = "NO";
    defparam add_4617_4.INJECT1_1 = "NO";
    CCU2D add_4617_2 (.A0(buf_r[1148]), .B0(buf_r[1177]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1149]), .B1(buf_r[1178]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62049), .S1(buf_x[1558]));
    defparam add_4617_2.INIT0 = 16'h7000;
    defparam add_4617_2.INIT1 = 16'h5666;
    defparam add_4617_2.INJECT1_0 = "NO";
    defparam add_4617_2.INJECT1_1 = "NO";
    CCU2D add_4616_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62047), 
          .S0(buf_x[1554]));
    defparam add_4616_cout.INIT0 = 16'h0000;
    defparam add_4616_cout.INIT1 = 16'h0000;
    defparam add_4616_cout.INJECT1_0 = "NO";
    defparam add_4616_cout.INJECT1_1 = "NO";
    CCU2D add_4616_30 (.A0(buf_r[1143]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_r[1144]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62046), .COUT(n62047), .S0(buf_x[1552]), .S1(buf_x[1553]));
    defparam add_4616_30.INIT0 = 16'hfaaa;
    defparam add_4616_30.INIT1 = 16'hfaaa;
    defparam add_4616_30.INJECT1_0 = "NO";
    defparam add_4616_30.INJECT1_1 = "NO";
    CCU2D add_4616_28 (.A0(buf_r[1112]), .B0(buf_r[1141]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1113]), .B1(buf_r[1142]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62045), .COUT(n62046), .S0(buf_x[1550]), 
          .S1(buf_x[1551]));
    defparam add_4616_28.INIT0 = 16'h5666;
    defparam add_4616_28.INIT1 = 16'h5666;
    defparam add_4616_28.INJECT1_0 = "NO";
    defparam add_4616_28.INJECT1_1 = "NO";
    CCU2D add_4616_26 (.A0(buf_r[1110]), .B0(buf_r[1139]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1111]), .B1(buf_r[1140]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62044), .COUT(n62045), .S0(buf_x[1548]), 
          .S1(buf_x[1549]));
    defparam add_4616_26.INIT0 = 16'h5666;
    defparam add_4616_26.INIT1 = 16'h5666;
    defparam add_4616_26.INJECT1_0 = "NO";
    defparam add_4616_26.INJECT1_1 = "NO";
    CCU2D add_4616_24 (.A0(buf_r[1108]), .B0(buf_r[1137]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1109]), .B1(buf_r[1138]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62043), .COUT(n62044), .S0(buf_x[1546]), 
          .S1(buf_x[1547]));
    defparam add_4616_24.INIT0 = 16'h5666;
    defparam add_4616_24.INIT1 = 16'h5666;
    defparam add_4616_24.INJECT1_0 = "NO";
    defparam add_4616_24.INJECT1_1 = "NO";
    CCU2D add_4616_22 (.A0(buf_r[1106]), .B0(buf_r[1135]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1107]), .B1(buf_r[1136]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62042), .COUT(n62043), .S0(buf_x[1544]), 
          .S1(buf_x[1545]));
    defparam add_4616_22.INIT0 = 16'h5666;
    defparam add_4616_22.INIT1 = 16'h5666;
    defparam add_4616_22.INJECT1_0 = "NO";
    defparam add_4616_22.INJECT1_1 = "NO";
    CCU2D add_4616_20 (.A0(buf_r[1104]), .B0(buf_r[1133]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1105]), .B1(buf_r[1134]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62041), .COUT(n62042), .S0(buf_x[1542]), 
          .S1(buf_x[1543]));
    defparam add_4616_20.INIT0 = 16'h5666;
    defparam add_4616_20.INIT1 = 16'h5666;
    defparam add_4616_20.INJECT1_0 = "NO";
    defparam add_4616_20.INJECT1_1 = "NO";
    CCU2D add_4616_18 (.A0(buf_r[1102]), .B0(buf_r[1131]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1103]), .B1(buf_r[1132]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62040), .COUT(n62041), .S0(buf_x[1540]), 
          .S1(buf_x[1541]));
    defparam add_4616_18.INIT0 = 16'h5666;
    defparam add_4616_18.INIT1 = 16'h5666;
    defparam add_4616_18.INJECT1_0 = "NO";
    defparam add_4616_18.INJECT1_1 = "NO";
    CCU2D add_4616_16 (.A0(buf_r[1100]), .B0(buf_r[1129]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1101]), .B1(buf_r[1130]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62039), .COUT(n62040), .S0(buf_x[1538]), 
          .S1(buf_x[1539]));
    defparam add_4616_16.INIT0 = 16'h5666;
    defparam add_4616_16.INIT1 = 16'h5666;
    defparam add_4616_16.INJECT1_0 = "NO";
    defparam add_4616_16.INJECT1_1 = "NO";
    CCU2D add_4616_14 (.A0(buf_r[1098]), .B0(buf_r[1127]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1099]), .B1(buf_r[1128]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62038), .COUT(n62039), .S0(buf_x[1536]), 
          .S1(buf_x[1537]));
    defparam add_4616_14.INIT0 = 16'h5666;
    defparam add_4616_14.INIT1 = 16'h5666;
    defparam add_4616_14.INJECT1_0 = "NO";
    defparam add_4616_14.INJECT1_1 = "NO";
    CCU2D add_4616_12 (.A0(buf_r[1096]), .B0(buf_r[1125]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1097]), .B1(buf_r[1126]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62037), .COUT(n62038), .S0(buf_x[1534]), 
          .S1(buf_x[1535]));
    defparam add_4616_12.INIT0 = 16'h5666;
    defparam add_4616_12.INIT1 = 16'h5666;
    defparam add_4616_12.INJECT1_0 = "NO";
    defparam add_4616_12.INJECT1_1 = "NO";
    CCU2D add_4616_10 (.A0(buf_r[1094]), .B0(buf_r[1123]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1095]), .B1(buf_r[1124]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62036), .COUT(n62037), .S0(buf_x[1532]), 
          .S1(buf_x[1533]));
    defparam add_4616_10.INIT0 = 16'h5666;
    defparam add_4616_10.INIT1 = 16'h5666;
    defparam add_4616_10.INJECT1_0 = "NO";
    defparam add_4616_10.INJECT1_1 = "NO";
    CCU2D add_4616_8 (.A0(buf_r[1092]), .B0(buf_r[1121]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1093]), .B1(buf_r[1122]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62035), .COUT(n62036), .S0(buf_x[1530]), 
          .S1(buf_x[1531]));
    defparam add_4616_8.INIT0 = 16'h5666;
    defparam add_4616_8.INIT1 = 16'h5666;
    defparam add_4616_8.INJECT1_0 = "NO";
    defparam add_4616_8.INJECT1_1 = "NO";
    CCU2D add_4616_6 (.A0(buf_r[1090]), .B0(buf_r[1119]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1091]), .B1(buf_r[1120]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62034), .COUT(n62035), .S0(buf_x[1528]), 
          .S1(buf_x[1529]));
    defparam add_4616_6.INIT0 = 16'h5666;
    defparam add_4616_6.INIT1 = 16'h5666;
    defparam add_4616_6.INJECT1_0 = "NO";
    defparam add_4616_6.INJECT1_1 = "NO";
    CCU2D add_4616_4 (.A0(buf_r[1088]), .B0(buf_r[1117]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1089]), .B1(buf_r[1118]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62033), .COUT(n62034), .S0(buf_x[1526]), 
          .S1(buf_x[1527]));
    defparam add_4616_4.INIT0 = 16'h5666;
    defparam add_4616_4.INIT1 = 16'h5666;
    defparam add_4616_4.INJECT1_0 = "NO";
    defparam add_4616_4.INJECT1_1 = "NO";
    CCU2D add_4616_2 (.A0(buf_r[1086]), .B0(buf_r[1115]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1087]), .B1(buf_r[1116]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62033), .S1(buf_x[1760]));
    defparam add_4616_2.INIT0 = 16'h7000;
    defparam add_4616_2.INIT1 = 16'h5666;
    defparam add_4616_2.INJECT1_0 = "NO";
    defparam add_4616_2.INJECT1_1 = "NO";
    CCU2D add_4615_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62031), 
          .S0(buf_x[1521]));
    defparam add_4615_cout.INIT0 = 16'h0000;
    defparam add_4615_cout.INIT1 = 16'h0000;
    defparam add_4615_cout.INJECT1_0 = "NO";
    defparam add_4615_cout.INJECT1_1 = "NO";
    CCU2D add_4615_30 (.A0(buf_r[1081]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_r[1082]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62030), .COUT(n62031), .S0(buf_x[1519]), .S1(buf_x[1520]));
    defparam add_4615_30.INIT0 = 16'hfaaa;
    defparam add_4615_30.INIT1 = 16'hfaaa;
    defparam add_4615_30.INJECT1_0 = "NO";
    defparam add_4615_30.INJECT1_1 = "NO";
    CCU2D add_4615_28 (.A0(buf_r[1050]), .B0(buf_r[1079]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1051]), .B1(buf_r[1080]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62029), .COUT(n62030), .S0(buf_x[1517]), 
          .S1(buf_x[1518]));
    defparam add_4615_28.INIT0 = 16'h5666;
    defparam add_4615_28.INIT1 = 16'h5666;
    defparam add_4615_28.INJECT1_0 = "NO";
    defparam add_4615_28.INJECT1_1 = "NO";
    CCU2D add_4615_26 (.A0(buf_r[1048]), .B0(buf_r[1077]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1049]), .B1(buf_r[1078]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62028), .COUT(n62029), .S0(buf_x[1515]), 
          .S1(buf_x[1516]));
    defparam add_4615_26.INIT0 = 16'h5666;
    defparam add_4615_26.INIT1 = 16'h5666;
    defparam add_4615_26.INJECT1_0 = "NO";
    defparam add_4615_26.INJECT1_1 = "NO";
    CCU2D add_4615_24 (.A0(buf_r[1046]), .B0(buf_r[1075]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1047]), .B1(buf_r[1076]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62027), .COUT(n62028), .S0(buf_x[1513]), 
          .S1(buf_x[1514]));
    defparam add_4615_24.INIT0 = 16'h5666;
    defparam add_4615_24.INIT1 = 16'h5666;
    defparam add_4615_24.INJECT1_0 = "NO";
    defparam add_4615_24.INJECT1_1 = "NO";
    CCU2D add_4615_22 (.A0(buf_r[1044]), .B0(buf_r[1073]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1045]), .B1(buf_r[1074]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62026), .COUT(n62027), .S0(buf_x[1511]), 
          .S1(buf_x[1512]));
    defparam add_4615_22.INIT0 = 16'h5666;
    defparam add_4615_22.INIT1 = 16'h5666;
    defparam add_4615_22.INJECT1_0 = "NO";
    defparam add_4615_22.INJECT1_1 = "NO";
    CCU2D add_4615_20 (.A0(buf_r[1042]), .B0(buf_r[1071]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1043]), .B1(buf_r[1072]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62025), .COUT(n62026), .S0(buf_x[1509]), 
          .S1(buf_x[1510]));
    defparam add_4615_20.INIT0 = 16'h5666;
    defparam add_4615_20.INIT1 = 16'h5666;
    defparam add_4615_20.INJECT1_0 = "NO";
    defparam add_4615_20.INJECT1_1 = "NO";
    CCU2D add_4615_18 (.A0(buf_r[1040]), .B0(buf_r[1069]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1041]), .B1(buf_r[1070]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62024), .COUT(n62025), .S0(buf_x[1507]), 
          .S1(buf_x[1508]));
    defparam add_4615_18.INIT0 = 16'h5666;
    defparam add_4615_18.INIT1 = 16'h5666;
    defparam add_4615_18.INJECT1_0 = "NO";
    defparam add_4615_18.INJECT1_1 = "NO";
    CCU2D add_4615_16 (.A0(buf_r[1038]), .B0(buf_r[1067]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1039]), .B1(buf_r[1068]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62023), .COUT(n62024), .S0(buf_x[1505]), 
          .S1(buf_x[1506]));
    defparam add_4615_16.INIT0 = 16'h5666;
    defparam add_4615_16.INIT1 = 16'h5666;
    defparam add_4615_16.INJECT1_0 = "NO";
    defparam add_4615_16.INJECT1_1 = "NO";
    CCU2D add_4615_14 (.A0(buf_r[1036]), .B0(buf_r[1065]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1037]), .B1(buf_r[1066]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62022), .COUT(n62023), .S0(buf_x[1503]), 
          .S1(buf_x[1504]));
    defparam add_4615_14.INIT0 = 16'h5666;
    defparam add_4615_14.INIT1 = 16'h5666;
    defparam add_4615_14.INJECT1_0 = "NO";
    defparam add_4615_14.INJECT1_1 = "NO";
    CCU2D add_4615_12 (.A0(buf_r[1034]), .B0(buf_r[1063]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1035]), .B1(buf_r[1064]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62021), .COUT(n62022), .S0(buf_x[1501]), 
          .S1(buf_x[1502]));
    defparam add_4615_12.INIT0 = 16'h5666;
    defparam add_4615_12.INIT1 = 16'h5666;
    defparam add_4615_12.INJECT1_0 = "NO";
    defparam add_4615_12.INJECT1_1 = "NO";
    CCU2D add_4615_10 (.A0(buf_r[1032]), .B0(buf_r[1061]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1033]), .B1(buf_r[1062]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62020), .COUT(n62021), .S0(buf_x[1499]), 
          .S1(buf_x[1500]));
    defparam add_4615_10.INIT0 = 16'h5666;
    defparam add_4615_10.INIT1 = 16'h5666;
    defparam add_4615_10.INJECT1_0 = "NO";
    defparam add_4615_10.INJECT1_1 = "NO";
    CCU2D add_4615_8 (.A0(buf_r[1030]), .B0(buf_r[1059]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1031]), .B1(buf_r[1060]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62019), .COUT(n62020), .S0(buf_x[1497]), 
          .S1(buf_x[1498]));
    defparam add_4615_8.INIT0 = 16'h5666;
    defparam add_4615_8.INIT1 = 16'h5666;
    defparam add_4615_8.INJECT1_0 = "NO";
    defparam add_4615_8.INJECT1_1 = "NO";
    CCU2D add_4615_6 (.A0(buf_r[1028]), .B0(buf_r[1057]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1029]), .B1(buf_r[1058]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62018), .COUT(n62019), .S0(buf_x[1495]), 
          .S1(buf_x[1496]));
    defparam add_4615_6.INIT0 = 16'h5666;
    defparam add_4615_6.INIT1 = 16'h5666;
    defparam add_4615_6.INJECT1_0 = "NO";
    defparam add_4615_6.INJECT1_1 = "NO";
    CCU2D add_4615_4 (.A0(buf_r[1026]), .B0(buf_r[1055]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1027]), .B1(buf_r[1056]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62017), .COUT(n62018), .S0(buf_x[1493]), 
          .S1(buf_x[1494]));
    defparam add_4615_4.INIT0 = 16'h5666;
    defparam add_4615_4.INIT1 = 16'h5666;
    defparam add_4615_4.INJECT1_0 = "NO";
    defparam add_4615_4.INJECT1_1 = "NO";
    CCU2D add_4615_2 (.A0(buf_r[1024]), .B0(buf_r[1053]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[1025]), .B1(buf_r[1054]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62017), .S1(buf_x[1492]));
    defparam add_4615_2.INIT0 = 16'h7000;
    defparam add_4615_2.INIT1 = 16'h5666;
    defparam add_4615_2.INJECT1_0 = "NO";
    defparam add_4615_2.INJECT1_1 = "NO";
    CCU2D add_4614_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62015), 
          .S0(buf_x[1488]));
    defparam add_4614_cout.INIT0 = 16'h0000;
    defparam add_4614_cout.INIT1 = 16'h0000;
    defparam add_4614_cout.INJECT1_0 = "NO";
    defparam add_4614_cout.INJECT1_1 = "NO";
    CCU2D add_4614_30 (.A0(buf_r[1019]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_r[1020]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62014), .COUT(n62015), .S0(buf_x[1486]), .S1(buf_x[1487]));
    defparam add_4614_30.INIT0 = 16'hfaaa;
    defparam add_4614_30.INIT1 = 16'hfaaa;
    defparam add_4614_30.INJECT1_0 = "NO";
    defparam add_4614_30.INJECT1_1 = "NO";
    CCU2D add_4614_28 (.A0(buf_r[988]), .B0(buf_r[1017]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[989]), .B1(buf_r[1018]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62013), .COUT(n62014), .S0(buf_x[1484]), 
          .S1(buf_x[1485]));
    defparam add_4614_28.INIT0 = 16'h5666;
    defparam add_4614_28.INIT1 = 16'h5666;
    defparam add_4614_28.INJECT1_0 = "NO";
    defparam add_4614_28.INJECT1_1 = "NO";
    CCU2D add_4614_26 (.A0(buf_r[986]), .B0(buf_r[1015]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[987]), .B1(buf_r[1016]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62012), .COUT(n62013), .S0(buf_x[1482]), 
          .S1(buf_x[1483]));
    defparam add_4614_26.INIT0 = 16'h5666;
    defparam add_4614_26.INIT1 = 16'h5666;
    defparam add_4614_26.INJECT1_0 = "NO";
    defparam add_4614_26.INJECT1_1 = "NO";
    CCU2D add_4614_24 (.A0(buf_r[984]), .B0(buf_r[1013]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[985]), .B1(buf_r[1014]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62011), .COUT(n62012), .S0(buf_x[1480]), 
          .S1(buf_x[1481]));
    defparam add_4614_24.INIT0 = 16'h5666;
    defparam add_4614_24.INIT1 = 16'h5666;
    defparam add_4614_24.INJECT1_0 = "NO";
    defparam add_4614_24.INJECT1_1 = "NO";
    CCU2D add_4614_22 (.A0(buf_r[982]), .B0(buf_r[1011]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[983]), .B1(buf_r[1012]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62010), .COUT(n62011), .S0(buf_x[1478]), 
          .S1(buf_x[1479]));
    defparam add_4614_22.INIT0 = 16'h5666;
    defparam add_4614_22.INIT1 = 16'h5666;
    defparam add_4614_22.INJECT1_0 = "NO";
    defparam add_4614_22.INJECT1_1 = "NO";
    CCU2D add_4614_20 (.A0(buf_r[980]), .B0(buf_r[1009]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[981]), .B1(buf_r[1010]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62009), .COUT(n62010), .S0(buf_x[1476]), 
          .S1(buf_x[1477]));
    defparam add_4614_20.INIT0 = 16'h5666;
    defparam add_4614_20.INIT1 = 16'h5666;
    defparam add_4614_20.INJECT1_0 = "NO";
    defparam add_4614_20.INJECT1_1 = "NO";
    CCU2D add_4614_18 (.A0(buf_r[978]), .B0(buf_r[1007]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[979]), .B1(buf_r[1008]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62008), .COUT(n62009), .S0(buf_x[1474]), 
          .S1(buf_x[1475]));
    defparam add_4614_18.INIT0 = 16'h5666;
    defparam add_4614_18.INIT1 = 16'h5666;
    defparam add_4614_18.INJECT1_0 = "NO";
    defparam add_4614_18.INJECT1_1 = "NO";
    CCU2D add_4614_16 (.A0(buf_r[976]), .B0(buf_r[1005]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[977]), .B1(buf_r[1006]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62007), .COUT(n62008), .S0(buf_x[1472]), 
          .S1(buf_x[1473]));
    defparam add_4614_16.INIT0 = 16'h5666;
    defparam add_4614_16.INIT1 = 16'h5666;
    defparam add_4614_16.INJECT1_0 = "NO";
    defparam add_4614_16.INJECT1_1 = "NO";
    CCU2D add_4614_14 (.A0(buf_r[974]), .B0(buf_r[1003]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[975]), .B1(buf_r[1004]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62006), .COUT(n62007), .S0(buf_x[1470]), 
          .S1(buf_x[1471]));
    defparam add_4614_14.INIT0 = 16'h5666;
    defparam add_4614_14.INIT1 = 16'h5666;
    defparam add_4614_14.INJECT1_0 = "NO";
    defparam add_4614_14.INJECT1_1 = "NO";
    CCU2D add_4614_12 (.A0(buf_r[972]), .B0(buf_r[1001]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[973]), .B1(buf_r[1002]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62005), .COUT(n62006), .S0(buf_x[1468]), 
          .S1(buf_x[1469]));
    defparam add_4614_12.INIT0 = 16'h5666;
    defparam add_4614_12.INIT1 = 16'h5666;
    defparam add_4614_12.INJECT1_0 = "NO";
    defparam add_4614_12.INJECT1_1 = "NO";
    CCU2D add_4614_10 (.A0(buf_r[970]), .B0(buf_r[999]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[971]), .B1(buf_r[1000]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62004), .COUT(n62005), .S0(buf_x[1466]), 
          .S1(buf_x[1467]));
    defparam add_4614_10.INIT0 = 16'h5666;
    defparam add_4614_10.INIT1 = 16'h5666;
    defparam add_4614_10.INJECT1_0 = "NO";
    defparam add_4614_10.INJECT1_1 = "NO";
    CCU2D add_4614_8 (.A0(buf_r[968]), .B0(buf_r[997]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[969]), .B1(buf_r[998]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62003), .COUT(n62004), .S0(buf_x[1464]), 
          .S1(buf_x[1465]));
    defparam add_4614_8.INIT0 = 16'h5666;
    defparam add_4614_8.INIT1 = 16'h5666;
    defparam add_4614_8.INJECT1_0 = "NO";
    defparam add_4614_8.INJECT1_1 = "NO";
    CCU2D add_4614_6 (.A0(buf_r[966]), .B0(buf_r[995]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[967]), .B1(buf_r[996]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62002), .COUT(n62003), .S0(buf_x[1462]), 
          .S1(buf_x[1463]));
    defparam add_4614_6.INIT0 = 16'h5666;
    defparam add_4614_6.INIT1 = 16'h5666;
    defparam add_4614_6.INJECT1_0 = "NO";
    defparam add_4614_6.INJECT1_1 = "NO";
    CCU2D add_4614_4 (.A0(buf_r[964]), .B0(buf_r[993]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[965]), .B1(buf_r[994]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62001), .COUT(n62002), .S0(buf_x[1460]), 
          .S1(buf_x[1461]));
    defparam add_4614_4.INIT0 = 16'h5666;
    defparam add_4614_4.INIT1 = 16'h5666;
    defparam add_4614_4.INJECT1_0 = "NO";
    defparam add_4614_4.INJECT1_1 = "NO";
    CCU2D add_4614_2 (.A0(buf_r[962]), .B0(buf_r[991]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[963]), .B1(buf_r[992]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62001));
    defparam add_4614_2.INIT0 = 16'h7000;
    defparam add_4614_2.INIT1 = 16'h5666;
    defparam add_4614_2.INJECT1_0 = "NO";
    defparam add_4614_2.INJECT1_1 = "NO";
    CCU2D add_4613_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[21]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62000), .S0(buf_x[1298]), .S1(buf_x[1299]));
    defparam add_4613_29.INIT0 = 16'h7888;
    defparam add_4613_29.INIT1 = 16'h0000;
    defparam add_4613_29.INJECT1_0 = "NO";
    defparam add_4613_29.INJECT1_1 = "NO";
    CCU2D add_4613_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[20]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[27]), .B1(nZ0_d2[20]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[21]), .CIN(n61999), .COUT(n62000), .S0(buf_x[1296]), 
          .S1(buf_x[1297]));
    defparam add_4613_27.INIT0 = 16'h7888;
    defparam add_4613_27.INIT1 = 16'h7888;
    defparam add_4613_27.INJECT1_0 = "NO";
    defparam add_4613_27.INJECT1_1 = "NO";
    CCU2D add_4613_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[20]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[25]), .B1(nZ0_d2[20]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[21]), .CIN(n61998), .COUT(n61999), .S0(buf_x[1294]), 
          .S1(buf_x[1295]));
    defparam add_4613_25.INIT0 = 16'h7888;
    defparam add_4613_25.INIT1 = 16'h7888;
    defparam add_4613_25.INJECT1_0 = "NO";
    defparam add_4613_25.INJECT1_1 = "NO";
    CCU2D add_4613_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[20]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[23]), .B1(nZ0_d2[20]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[21]), .CIN(n61997), .COUT(n61998), .S0(buf_x[1292]), 
          .S1(buf_x[1293]));
    defparam add_4613_23.INIT0 = 16'h7888;
    defparam add_4613_23.INIT1 = 16'h7888;
    defparam add_4613_23.INJECT1_0 = "NO";
    defparam add_4613_23.INJECT1_1 = "NO";
    CCU2D add_4613_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[20]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[21]), .B1(nZ0_d2[20]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[21]), .CIN(n61996), .COUT(n61997), .S0(buf_x[1290]), 
          .S1(buf_x[1291]));
    defparam add_4613_21.INIT0 = 16'h7888;
    defparam add_4613_21.INIT1 = 16'h7888;
    defparam add_4613_21.INJECT1_0 = "NO";
    defparam add_4613_21.INJECT1_1 = "NO";
    CCU2D add_4613_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[20]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[19]), .B1(nZ0_d2[20]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[21]), .CIN(n61995), .COUT(n61996), .S0(buf_x[1288]), 
          .S1(buf_x[1289]));
    defparam add_4613_19.INIT0 = 16'h7888;
    defparam add_4613_19.INIT1 = 16'h7888;
    defparam add_4613_19.INJECT1_0 = "NO";
    defparam add_4613_19.INJECT1_1 = "NO";
    CCU2D add_4613_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[20]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[17]), .B1(nZ0_d2[20]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[21]), .CIN(n61994), .COUT(n61995), .S0(buf_x[1286]), 
          .S1(buf_x[1287]));
    defparam add_4613_17.INIT0 = 16'h7888;
    defparam add_4613_17.INIT1 = 16'h7888;
    defparam add_4613_17.INJECT1_0 = "NO";
    defparam add_4613_17.INJECT1_1 = "NO";
    CCU2D add_4613_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[20]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[15]), .B1(nZ0_d2[20]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[21]), .CIN(n61993), .COUT(n61994), .S0(buf_x[1284]), 
          .S1(buf_x[1285]));
    defparam add_4613_15.INIT0 = 16'h7888;
    defparam add_4613_15.INIT1 = 16'h7888;
    defparam add_4613_15.INJECT1_0 = "NO";
    defparam add_4613_15.INJECT1_1 = "NO";
    CCU2D add_4613_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[20]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[13]), .B1(nZ0_d2[20]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[21]), .CIN(n61992), .COUT(n61993), .S0(buf_x[1282]), 
          .S1(buf_x[1283]));
    defparam add_4613_13.INIT0 = 16'h7888;
    defparam add_4613_13.INIT1 = 16'h7888;
    defparam add_4613_13.INJECT1_0 = "NO";
    defparam add_4613_13.INJECT1_1 = "NO";
    CCU2D add_4613_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[20]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[11]), .B1(nZ0_d2[20]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[21]), .CIN(n61991), .COUT(n61992), .S0(buf_x[1280]), 
          .S1(buf_x[1281]));
    defparam add_4613_11.INIT0 = 16'h7888;
    defparam add_4613_11.INIT1 = 16'h7888;
    defparam add_4613_11.INJECT1_0 = "NO";
    defparam add_4613_11.INJECT1_1 = "NO";
    CCU2D add_4613_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[20]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[9]), .B1(nZ0_d2[20]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[21]), .CIN(n61990), .COUT(n61991), .S0(buf_x[1278]), 
          .S1(buf_x[1279]));
    defparam add_4613_9.INIT0 = 16'h7888;
    defparam add_4613_9.INIT1 = 16'h7888;
    defparam add_4613_9.INJECT1_0 = "NO";
    defparam add_4613_9.INJECT1_1 = "NO";
    CCU2D add_4613_7 (.A0(nEY1_d2[6]), .B0(nZ0_d2[20]), .C0(nEY1_d2[5]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[7]), .B1(nZ0_d2[20]), .C1(nEY1_d2[6]), 
          .D1(nZ0_d2[21]), .CIN(n61989), .COUT(n61990), .S0(buf_x[1276]), 
          .S1(buf_x[1277]));
    defparam add_4613_7.INIT0 = 16'h7888;
    defparam add_4613_7.INIT1 = 16'h7888;
    defparam add_4613_7.INJECT1_0 = "NO";
    defparam add_4613_7.INJECT1_1 = "NO";
    CCU2D add_4613_5 (.A0(nEY1_d2[4]), .B0(nZ0_d2[20]), .C0(nEY1_d2[3]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[5]), .B1(nZ0_d2[20]), .C1(nEY1_d2[4]), 
          .D1(nZ0_d2[21]), .CIN(n61988), .COUT(n61989), .S0(buf_x[1274]), 
          .S1(buf_x[1275]));
    defparam add_4613_5.INIT0 = 16'h7888;
    defparam add_4613_5.INIT1 = 16'h7888;
    defparam add_4613_5.INJECT1_0 = "NO";
    defparam add_4613_5.INJECT1_1 = "NO";
    CCU2D add_4613_3 (.A0(nEY1_d2[2]), .B0(nZ0_d2[20]), .C0(nEY1_d2[1]), 
          .D0(nZ0_d2[21]), .A1(nEY1_d2[3]), .B1(nZ0_d2[20]), .C1(nEY1_d2[2]), 
          .D1(nZ0_d2[21]), .CIN(n61987), .COUT(n61988), .S0(buf_x[1272]), 
          .S1(buf_x[1273]));
    defparam add_4613_3.INIT0 = 16'h7888;
    defparam add_4613_3.INIT1 = 16'h7888;
    defparam add_4613_3.INJECT1_0 = "NO";
    defparam add_4613_3.INJECT1_1 = "NO";
    CCU2D add_4613_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(nEY1_d2[1]), .B1(nZ0_d2[20]), .C1(nEY1_d2[0]), .D1(nZ0_d2[21]), 
          .COUT(n61987), .S1(buf_x[1271]));
    defparam add_4613_1.INIT0 = 16'hF000;
    defparam add_4613_1.INIT1 = 16'h7888;
    defparam add_4613_1.INJECT1_0 = "NO";
    defparam add_4613_1.INJECT1_1 = "NO";
    CCU2D add_4612_29 (.A0(nEY1_d2[27]), .B0(nZ0_d2[19]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61986), .S0(buf_x[1267]), .S1(buf_x[1268]));
    defparam add_4612_29.INIT0 = 16'h7888;
    defparam add_4612_29.INIT1 = 16'h0000;
    defparam add_4612_29.INJECT1_0 = "NO";
    defparam add_4612_29.INJECT1_1 = "NO";
    CCU2D add_4612_27 (.A0(nEY1_d2[26]), .B0(nZ0_d2[18]), .C0(nEY1_d2[25]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[27]), .B1(nZ0_d2[18]), .C1(nEY1_d2[26]), 
          .D1(nZ0_d2[19]), .CIN(n61985), .COUT(n61986), .S0(buf_x[1265]), 
          .S1(buf_x[1266]));
    defparam add_4612_27.INIT0 = 16'h7888;
    defparam add_4612_27.INIT1 = 16'h7888;
    defparam add_4612_27.INJECT1_0 = "NO";
    defparam add_4612_27.INJECT1_1 = "NO";
    CCU2D add_4612_25 (.A0(nEY1_d2[24]), .B0(nZ0_d2[18]), .C0(nEY1_d2[23]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[25]), .B1(nZ0_d2[18]), .C1(nEY1_d2[24]), 
          .D1(nZ0_d2[19]), .CIN(n61984), .COUT(n61985), .S0(buf_x[1263]), 
          .S1(buf_x[1264]));
    defparam add_4612_25.INIT0 = 16'h7888;
    defparam add_4612_25.INIT1 = 16'h7888;
    defparam add_4612_25.INJECT1_0 = "NO";
    defparam add_4612_25.INJECT1_1 = "NO";
    CCU2D add_4612_23 (.A0(nEY1_d2[22]), .B0(nZ0_d2[18]), .C0(nEY1_d2[21]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[23]), .B1(nZ0_d2[18]), .C1(nEY1_d2[22]), 
          .D1(nZ0_d2[19]), .CIN(n61983), .COUT(n61984), .S0(buf_x[1261]), 
          .S1(buf_x[1262]));
    defparam add_4612_23.INIT0 = 16'h7888;
    defparam add_4612_23.INIT1 = 16'h7888;
    defparam add_4612_23.INJECT1_0 = "NO";
    defparam add_4612_23.INJECT1_1 = "NO";
    CCU2D add_4612_21 (.A0(nEY1_d2[20]), .B0(nZ0_d2[18]), .C0(nEY1_d2[19]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[21]), .B1(nZ0_d2[18]), .C1(nEY1_d2[20]), 
          .D1(nZ0_d2[19]), .CIN(n61982), .COUT(n61983), .S0(buf_x[1259]), 
          .S1(buf_x[1260]));
    defparam add_4612_21.INIT0 = 16'h7888;
    defparam add_4612_21.INIT1 = 16'h7888;
    defparam add_4612_21.INJECT1_0 = "NO";
    defparam add_4612_21.INJECT1_1 = "NO";
    CCU2D add_4612_19 (.A0(nEY1_d2[18]), .B0(nZ0_d2[18]), .C0(nEY1_d2[17]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[19]), .B1(nZ0_d2[18]), .C1(nEY1_d2[18]), 
          .D1(nZ0_d2[19]), .CIN(n61981), .COUT(n61982), .S0(buf_x[1257]), 
          .S1(buf_x[1258]));
    defparam add_4612_19.INIT0 = 16'h7888;
    defparam add_4612_19.INIT1 = 16'h7888;
    defparam add_4612_19.INJECT1_0 = "NO";
    defparam add_4612_19.INJECT1_1 = "NO";
    CCU2D add_4612_17 (.A0(nEY1_d2[16]), .B0(nZ0_d2[18]), .C0(nEY1_d2[15]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[17]), .B1(nZ0_d2[18]), .C1(nEY1_d2[16]), 
          .D1(nZ0_d2[19]), .CIN(n61980), .COUT(n61981), .S0(buf_x[1255]), 
          .S1(buf_x[1256]));
    defparam add_4612_17.INIT0 = 16'h7888;
    defparam add_4612_17.INIT1 = 16'h7888;
    defparam add_4612_17.INJECT1_0 = "NO";
    defparam add_4612_17.INJECT1_1 = "NO";
    CCU2D add_4612_15 (.A0(nEY1_d2[14]), .B0(nZ0_d2[18]), .C0(nEY1_d2[13]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[15]), .B1(nZ0_d2[18]), .C1(nEY1_d2[14]), 
          .D1(nZ0_d2[19]), .CIN(n61979), .COUT(n61980), .S0(buf_x[1253]), 
          .S1(buf_x[1254]));
    defparam add_4612_15.INIT0 = 16'h7888;
    defparam add_4612_15.INIT1 = 16'h7888;
    defparam add_4612_15.INJECT1_0 = "NO";
    defparam add_4612_15.INJECT1_1 = "NO";
    CCU2D add_4612_13 (.A0(nEY1_d2[12]), .B0(nZ0_d2[18]), .C0(nEY1_d2[11]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[13]), .B1(nZ0_d2[18]), .C1(nEY1_d2[12]), 
          .D1(nZ0_d2[19]), .CIN(n61978), .COUT(n61979), .S0(buf_x[1251]), 
          .S1(buf_x[1252]));
    defparam add_4612_13.INIT0 = 16'h7888;
    defparam add_4612_13.INIT1 = 16'h7888;
    defparam add_4612_13.INJECT1_0 = "NO";
    defparam add_4612_13.INJECT1_1 = "NO";
    CCU2D add_4612_11 (.A0(nEY1_d2[10]), .B0(nZ0_d2[18]), .C0(nEY1_d2[9]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[11]), .B1(nZ0_d2[18]), .C1(nEY1_d2[10]), 
          .D1(nZ0_d2[19]), .CIN(n61977), .COUT(n61978), .S0(buf_x[1249]), 
          .S1(buf_x[1250]));
    defparam add_4612_11.INIT0 = 16'h7888;
    defparam add_4612_11.INIT1 = 16'h7888;
    defparam add_4612_11.INJECT1_0 = "NO";
    defparam add_4612_11.INJECT1_1 = "NO";
    CCU2D add_4612_9 (.A0(nEY1_d2[8]), .B0(nZ0_d2[18]), .C0(nEY1_d2[7]), 
          .D0(nZ0_d2[19]), .A1(nEY1_d2[9]), .B1(nZ0_d2[18]), .C1(nEY1_d2[8]), 
          .D1(nZ0_d2[19]), .CIN(n61976), .COUT(n61977), .S0(buf_x[1247]), 
          .S1(buf_x[1248]));
    defparam add_4612_9.INIT0 = 16'h7888;
    defparam add_4612_9.INIT1 = 16'h7888;
    defparam add_4612_9.INJECT1_0 = "NO";
    defparam add_4612_9.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \mult_clk(9,35,true,false,-1,2) 
//

module \mult_clk(9,35,true,false,-1,2)  (\buf_x[623] , clock, nK_b0, GND_net, 
            \nKLog2_c0[34] , \nKLog2_c0[32] , \nKLog2_c0[33] , \nKLog2_c0[30] , 
            \nKLog2_c0[31] , \nKLog2_c0[28] , \nKLog2_c0[29] , \nKLog2_c0[26] , 
            \nKLog2_c0[27] , \nKLog2_c0[24] , \nKLog2_c0[25] , \nKLog2_c0[22] , 
            \nKLog2_c0[23] , \nKLog2_c0[20] , \nKLog2_c0[21] , \nKLog2_c0[18] , 
            \nKLog2_c0[19] , \nKLog2_c0[16] , \nKLog2_c0[17] , \nKLog2_c0[14] , 
            \nKLog2_c0[15] , \nKLog2_c0[12] , \nKLog2_c0[13] , \nKLog2_c0[10] , 
            \nKLog2_c0[11] , \nKLog2_c0[9] , \buf_x[699] , \buf_x[689] , 
            \buf_x[737] , \buf_x[727] , \buf_x[651] , \buf_x[661] , 
            \buf_x[613] , \nKLog2_c0[7] , \buf_r[936] , \nKLog2_c0[8] );
    output \buf_x[623] ;
    input clock;
    input [8:0]nK_b0;
    input GND_net;
    output \nKLog2_c0[34] ;
    output \nKLog2_c0[32] ;
    output \nKLog2_c0[33] ;
    output \nKLog2_c0[30] ;
    output \nKLog2_c0[31] ;
    output \nKLog2_c0[28] ;
    output \nKLog2_c0[29] ;
    output \nKLog2_c0[26] ;
    output \nKLog2_c0[27] ;
    output \nKLog2_c0[24] ;
    output \nKLog2_c0[25] ;
    output \nKLog2_c0[22] ;
    output \nKLog2_c0[23] ;
    output \nKLog2_c0[20] ;
    output \nKLog2_c0[21] ;
    output \nKLog2_c0[18] ;
    output \nKLog2_c0[19] ;
    output \nKLog2_c0[16] ;
    output \nKLog2_c0[17] ;
    output \nKLog2_c0[14] ;
    output \nKLog2_c0[15] ;
    output \nKLog2_c0[12] ;
    output \nKLog2_c0[13] ;
    output \nKLog2_c0[10] ;
    output \nKLog2_c0[11] ;
    output \nKLog2_c0[9] ;
    output \buf_x[699] ;
    output \buf_x[689] ;
    output \buf_x[737] ;
    output \buf_x[727] ;
    output \buf_x[651] ;
    output \buf_x[661] ;
    output \buf_x[613] ;
    output \nKLog2_c0[7] ;
    input \buf_r[936] ;
    output \nKLog2_c0[8] ;
    
    wire [1195:0]buf_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [1195:0]buf_r;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(337[10:15])
    
    wire n62543, n62542, n62541, n62540, n62539, n62538, n62537, 
        n62536, n62535, n62534, n62533, n62532, n62531, n61825, 
        n61824, n61823, n61822, n61821, n61820, n61819, n61818, 
        n61817, n61816, n61815, n61814, n61813, n61812, n61811, 
        n61809, n61808, n61807, n61806, n61805, n61804, n61803, 
        n61802, n61801, n61800, n61799, n61798, n61797, n61794, 
        n61793, n61792, n61791, n61790, n61789, n61788, n61787, 
        n61786, n61785, n61784, n61783, n61782, n61781, n61780, 
        n61764, n61763, n61762, n61761, n61760, n61759, n61758, 
        n61757, n61756, n61749, n61748, n61747, n61746, n61745, 
        n61744, n61743, n61742, n61741, n61740, n61739, n61707, 
        n61706, n61705, n61704, n61703, n61702, n61701, n61700, 
        n61699, n61698, n61697, n61696, n61498, n61497, n61496, 
        n61495, n61494, n61493, n61492, n61491, n61490, n61489;
    
    FD1S3AX nK_b1_i1 (.D(nK_b0[0]), .CK(clock), .Q(\buf_x[623] ));
    defparam nK_b1_i1.GSR = "DISABLED";
    FD1S3AX buf_r_976__183 (.D(buf_x[1002]), .CK(clock), .Q(buf_x[1100]));
    defparam buf_r_976__183.GSR = "DISABLED";
    FD1S3AX buf_r_966__193 (.D(buf_x[966]), .CK(clock), .Q(buf_r[966]));
    defparam buf_r_966__193.GSR = "DISABLED";
    FD1S3AX buf_r_965__194 (.D(buf_x[965]), .CK(clock), .Q(buf_r[965]));
    defparam buf_r_965__194.GSR = "DISABLED";
    FD1S3AX buf_r_964__195 (.D(buf_x[964]), .CK(clock), .Q(buf_r[964]));
    defparam buf_r_964__195.GSR = "DISABLED";
    FD1S3AX buf_r_963__196 (.D(buf_x[963]), .CK(clock), .Q(buf_r[963]));
    defparam buf_r_963__196.GSR = "DISABLED";
    FD1S3AX buf_r_962__197 (.D(buf_x[962]), .CK(clock), .Q(buf_r[962]));
    defparam buf_r_962__197.GSR = "DISABLED";
    FD1S3AX buf_r_961__198 (.D(buf_x[961]), .CK(clock), .Q(buf_r[961]));
    defparam buf_r_961__198.GSR = "DISABLED";
    FD1S3AX buf_r_960__199 (.D(buf_x[960]), .CK(clock), .Q(buf_r[960]));
    defparam buf_r_960__199.GSR = "DISABLED";
    FD1S3AX buf_r_959__200 (.D(buf_x[959]), .CK(clock), .Q(buf_r[959]));
    defparam buf_r_959__200.GSR = "DISABLED";
    FD1S3AX buf_r_958__201 (.D(buf_x[958]), .CK(clock), .Q(buf_r[958]));
    defparam buf_r_958__201.GSR = "DISABLED";
    FD1S3AX buf_r_957__202 (.D(buf_x[957]), .CK(clock), .Q(buf_r[957]));
    defparam buf_r_957__202.GSR = "DISABLED";
    FD1S3AX buf_r_956__203 (.D(buf_x[956]), .CK(clock), .Q(buf_r[956]));
    defparam buf_r_956__203.GSR = "DISABLED";
    FD1S3AX buf_r_955__204 (.D(buf_x[955]), .CK(clock), .Q(buf_r[955]));
    defparam buf_r_955__204.GSR = "DISABLED";
    FD1S3AX buf_r_954__205 (.D(buf_x[954]), .CK(clock), .Q(buf_r[954]));
    defparam buf_r_954__205.GSR = "DISABLED";
    FD1S3AX buf_r_953__206 (.D(buf_x[953]), .CK(clock), .Q(buf_r[953]));
    defparam buf_r_953__206.GSR = "DISABLED";
    FD1S3AX buf_r_952__207 (.D(buf_x[952]), .CK(clock), .Q(buf_r[952]));
    defparam buf_r_952__207.GSR = "DISABLED";
    FD1S3AX buf_r_951__208 (.D(buf_x[951]), .CK(clock), .Q(buf_r[951]));
    defparam buf_r_951__208.GSR = "DISABLED";
    FD1S3AX buf_r_950__209 (.D(buf_x[950]), .CK(clock), .Q(buf_r[950]));
    defparam buf_r_950__209.GSR = "DISABLED";
    FD1S3AX buf_r_949__210 (.D(buf_x[948]), .CK(clock), .Q(buf_r[949]));
    defparam buf_r_949__210.GSR = "DISABLED";
    FD1S3AX buf_r_947__212 (.D(buf_x[947]), .CK(clock), .Q(buf_r[947]));
    defparam buf_r_947__212.GSR = "DISABLED";
    FD1S3AX buf_r_946__213 (.D(buf_x[946]), .CK(clock), .Q(buf_r[946]));
    defparam buf_r_946__213.GSR = "DISABLED";
    FD1S3AX buf_r_945__214 (.D(buf_x[945]), .CK(clock), .Q(buf_r[945]));
    defparam buf_r_945__214.GSR = "DISABLED";
    FD1S3AX buf_r_944__215 (.D(buf_x[944]), .CK(clock), .Q(buf_r[944]));
    defparam buf_r_944__215.GSR = "DISABLED";
    FD1S3AX buf_r_943__216 (.D(buf_x[943]), .CK(clock), .Q(buf_r[943]));
    defparam buf_r_943__216.GSR = "DISABLED";
    FD1S3AX buf_r_942__217 (.D(buf_x[942]), .CK(clock), .Q(buf_r[942]));
    defparam buf_r_942__217.GSR = "DISABLED";
    FD1S3AX buf_r_941__218 (.D(buf_x[941]), .CK(clock), .Q(buf_r[941]));
    defparam buf_r_941__218.GSR = "DISABLED";
    FD1S3AX buf_r_940__219 (.D(buf_x[940]), .CK(clock), .Q(buf_r[940]));
    defparam buf_r_940__219.GSR = "DISABLED";
    FD1S3AX buf_r_939__220 (.D(buf_x[939]), .CK(clock), .Q(buf_r[939]));
    defparam buf_r_939__220.GSR = "DISABLED";
    FD1S3AX buf_r_938__221 (.D(buf_x[938]), .CK(clock), .Q(buf_r[938]));
    defparam buf_r_938__221.GSR = "DISABLED";
    FD1S3AX buf_r_937__222 (.D(buf_x[937]), .CK(clock), .Q(buf_r[937]));
    defparam buf_r_937__222.GSR = "DISABLED";
    FD1S3AX buf_r_930__229 (.D(buf_x[930]), .CK(clock), .Q(buf_r[930]));
    defparam buf_r_930__229.GSR = "DISABLED";
    FD1S3AX buf_r_929__230 (.D(buf_x[929]), .CK(clock), .Q(buf_r[929]));
    defparam buf_r_929__230.GSR = "DISABLED";
    FD1S3AX buf_r_928__231 (.D(buf_x[928]), .CK(clock), .Q(buf_r[928]));
    defparam buf_r_928__231.GSR = "DISABLED";
    FD1S3AX buf_r_927__232 (.D(buf_x[927]), .CK(clock), .Q(buf_r[927]));
    defparam buf_r_927__232.GSR = "DISABLED";
    FD1S3AX buf_r_926__233 (.D(buf_x[926]), .CK(clock), .Q(buf_r[926]));
    defparam buf_r_926__233.GSR = "DISABLED";
    FD1S3AX buf_r_925__234 (.D(buf_x[925]), .CK(clock), .Q(buf_r[925]));
    defparam buf_r_925__234.GSR = "DISABLED";
    FD1S3AX buf_r_924__235 (.D(buf_x[924]), .CK(clock), .Q(buf_r[924]));
    defparam buf_r_924__235.GSR = "DISABLED";
    FD1S3AX buf_r_923__236 (.D(buf_x[923]), .CK(clock), .Q(buf_r[923]));
    defparam buf_r_923__236.GSR = "DISABLED";
    FD1S3AX buf_r_922__237 (.D(buf_x[922]), .CK(clock), .Q(buf_r[922]));
    defparam buf_r_922__237.GSR = "DISABLED";
    FD1S3AX buf_r_921__238 (.D(buf_x[921]), .CK(clock), .Q(buf_r[921]));
    defparam buf_r_921__238.GSR = "DISABLED";
    FD1S3AX buf_r_920__239 (.D(buf_x[920]), .CK(clock), .Q(buf_r[920]));
    defparam buf_r_920__239.GSR = "DISABLED";
    FD1S3AX buf_r_919__240 (.D(buf_x[919]), .CK(clock), .Q(buf_r[919]));
    defparam buf_r_919__240.GSR = "DISABLED";
    FD1S3AX buf_r_918__241 (.D(buf_x[918]), .CK(clock), .Q(buf_r[918]));
    defparam buf_r_918__241.GSR = "DISABLED";
    FD1S3AX buf_r_917__242 (.D(buf_x[917]), .CK(clock), .Q(buf_r[917]));
    defparam buf_r_917__242.GSR = "DISABLED";
    FD1S3AX buf_r_916__243 (.D(buf_x[916]), .CK(clock), .Q(buf_r[916]));
    defparam buf_r_916__243.GSR = "DISABLED";
    FD1S3AX buf_r_915__244 (.D(buf_x[915]), .CK(clock), .Q(buf_r[915]));
    defparam buf_r_915__244.GSR = "DISABLED";
    FD1S3AX buf_r_914__245 (.D(buf_x[914]), .CK(clock), .Q(buf_r[914]));
    defparam buf_r_914__245.GSR = "DISABLED";
    FD1S3AX buf_r_913__246 (.D(buf_x[913]), .CK(clock), .Q(buf_r[913]));
    defparam buf_r_913__246.GSR = "DISABLED";
    FD1S3AX buf_r_912__247 (.D(buf_x[912]), .CK(clock), .Q(buf_r[912]));
    defparam buf_r_912__247.GSR = "DISABLED";
    FD1S3AX buf_r_911__248 (.D(buf_x[911]), .CK(clock), .Q(buf_r[911]));
    defparam buf_r_911__248.GSR = "DISABLED";
    FD1S3AX buf_r_910__249 (.D(buf_x[910]), .CK(clock), .Q(buf_r[910]));
    defparam buf_r_910__249.GSR = "DISABLED";
    FD1S3AX buf_r_909__250 (.D(buf_x[908]), .CK(clock), .Q(buf_r[909]));
    defparam buf_r_909__250.GSR = "DISABLED";
    FD1S3AX buf_r_907__252 (.D(buf_x[907]), .CK(clock), .Q(buf_r[907]));
    defparam buf_r_907__252.GSR = "DISABLED";
    FD1S3AX buf_r_906__253 (.D(buf_x[906]), .CK(clock), .Q(buf_r[906]));
    defparam buf_r_906__253.GSR = "DISABLED";
    FD1S3AX buf_r_905__254 (.D(buf_x[905]), .CK(clock), .Q(buf_r[905]));
    defparam buf_r_905__254.GSR = "DISABLED";
    FD1S3AX buf_r_904__255 (.D(buf_x[904]), .CK(clock), .Q(buf_r[904]));
    defparam buf_r_904__255.GSR = "DISABLED";
    FD1S3AX buf_r_903__256 (.D(buf_x[903]), .CK(clock), .Q(buf_r[903]));
    defparam buf_r_903__256.GSR = "DISABLED";
    FD1S3AX buf_r_902__257 (.D(buf_x[902]), .CK(clock), .Q(buf_r[902]));
    defparam buf_r_902__257.GSR = "DISABLED";
    FD1S3AX buf_r_901__258 (.D(buf_x[901]), .CK(clock), .Q(buf_r[901]));
    defparam buf_r_901__258.GSR = "DISABLED";
    FD1S3AX buf_r_900__259 (.D(buf_x[900]), .CK(clock), .Q(buf_r[900]));
    defparam buf_r_900__259.GSR = "DISABLED";
    CCU2D add_4626_28 (.A0(buf_x[1090]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62543), .S0(\nKLog2_c0[34] ));
    defparam add_4626_28.INIT0 = 16'h5666;
    defparam add_4626_28.INIT1 = 16'h0000;
    defparam add_4626_28.INJECT1_0 = "NO";
    defparam add_4626_28.INJECT1_1 = "NO";
    CCU2D add_4626_26 (.A0(buf_x[1088]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1089]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62542), .COUT(n62543), .S0(\nKLog2_c0[32] ), .S1(\nKLog2_c0[33] ));
    defparam add_4626_26.INIT0 = 16'h5aaa;
    defparam add_4626_26.INIT1 = 16'h5aaa;
    defparam add_4626_26.INJECT1_0 = "NO";
    defparam add_4626_26.INJECT1_1 = "NO";
    CCU2D add_4626_24 (.A0(buf_x[1086]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1087]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62541), .COUT(n62542), .S0(\nKLog2_c0[30] ), 
          .S1(\nKLog2_c0[31] ));
    defparam add_4626_24.INIT0 = 16'h5666;
    defparam add_4626_24.INIT1 = 16'h5aaa;
    defparam add_4626_24.INJECT1_0 = "NO";
    defparam add_4626_24.INJECT1_1 = "NO";
    CCU2D add_4626_22 (.A0(buf_x[1084]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1085]), .B1(buf_x[1100]), .C1(GND_net), .D1(GND_net), 
          .CIN(n62540), .COUT(n62541), .S0(\nKLog2_c0[28] ), .S1(\nKLog2_c0[29] ));
    defparam add_4626_22.INIT0 = 16'h5aaa;
    defparam add_4626_22.INIT1 = 16'h5666;
    defparam add_4626_22.INJECT1_0 = "NO";
    defparam add_4626_22.INJECT1_1 = "NO";
    CCU2D add_4626_20 (.A0(buf_x[1082]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1083]), .B1(buf_x[1100]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62539), .COUT(n62540), .S0(\nKLog2_c0[26] ), 
          .S1(\nKLog2_c0[27] ));
    defparam add_4626_20.INIT0 = 16'h5666;
    defparam add_4626_20.INIT1 = 16'h5666;
    defparam add_4626_20.INJECT1_0 = "NO";
    defparam add_4626_20.INJECT1_1 = "NO";
    CCU2D add_4626_18 (.A0(buf_x[1080]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1081]), .B1(buf_x[1100]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62538), .COUT(n62539), .S0(\nKLog2_c0[24] ), 
          .S1(\nKLog2_c0[25] ));
    defparam add_4626_18.INIT0 = 16'h5666;
    defparam add_4626_18.INIT1 = 16'h5666;
    defparam add_4626_18.INJECT1_0 = "NO";
    defparam add_4626_18.INJECT1_1 = "NO";
    CCU2D add_4626_16 (.A0(buf_x[1078]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1079]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62537), .COUT(n62538), .S0(\nKLog2_c0[22] ), 
          .S1(\nKLog2_c0[23] ));
    defparam add_4626_16.INIT0 = 16'h5666;
    defparam add_4626_16.INIT1 = 16'h5aaa;
    defparam add_4626_16.INJECT1_0 = "NO";
    defparam add_4626_16.INJECT1_1 = "NO";
    CCU2D add_4626_14 (.A0(buf_x[1076]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1077]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62536), .COUT(n62537), .S0(\nKLog2_c0[20] ), .S1(\nKLog2_c0[21] ));
    defparam add_4626_14.INIT0 = 16'h5aaa;
    defparam add_4626_14.INIT1 = 16'h5aaa;
    defparam add_4626_14.INJECT1_0 = "NO";
    defparam add_4626_14.INJECT1_1 = "NO";
    CCU2D add_4626_12 (.A0(buf_x[1074]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1075]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62535), .COUT(n62536), .S0(\nKLog2_c0[18] ), .S1(\nKLog2_c0[19] ));
    defparam add_4626_12.INIT0 = 16'h5aaa;
    defparam add_4626_12.INIT1 = 16'h5aaa;
    defparam add_4626_12.INJECT1_0 = "NO";
    defparam add_4626_12.INJECT1_1 = "NO";
    CCU2D add_4626_10 (.A0(buf_x[1072]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1073]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62534), .COUT(n62535), .S0(\nKLog2_c0[16] ), .S1(\nKLog2_c0[17] ));
    defparam add_4626_10.INIT0 = 16'h5aaa;
    defparam add_4626_10.INIT1 = 16'h5aaa;
    defparam add_4626_10.INJECT1_0 = "NO";
    defparam add_4626_10.INJECT1_1 = "NO";
    CCU2D add_4626_8 (.A0(buf_x[1070]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1071]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62533), .COUT(n62534), .S0(\nKLog2_c0[14] ), 
          .S1(\nKLog2_c0[15] ));
    defparam add_4626_8.INIT0 = 16'h5666;
    defparam add_4626_8.INIT1 = 16'h5aaa;
    defparam add_4626_8.INJECT1_0 = "NO";
    defparam add_4626_8.INJECT1_1 = "NO";
    CCU2D add_4626_6 (.A0(buf_x[1068]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1069]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62532), .COUT(n62533), .S0(\nKLog2_c0[12] ), .S1(\nKLog2_c0[13] ));
    defparam add_4626_6.INIT0 = 16'h5aaa;
    defparam add_4626_6.INIT1 = 16'h5aaa;
    defparam add_4626_6.INJECT1_0 = "NO";
    defparam add_4626_6.INJECT1_1 = "NO";
    CCU2D add_4626_4 (.A0(buf_x[1066]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[1067]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62531), .COUT(n62532), .S0(\nKLog2_c0[10] ), .S1(\nKLog2_c0[11] ));
    defparam add_4626_4.INIT0 = 16'h5aaa;
    defparam add_4626_4.INIT1 = 16'h5aaa;
    defparam add_4626_4.INJECT1_0 = "NO";
    defparam add_4626_4.INJECT1_1 = "NO";
    CCU2D add_4626_2 (.A0(buf_x[1064]), .B0(buf_x[1100]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[1065]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n62531), .S1(\nKLog2_c0[9] ));
    defparam add_4626_2.INIT0 = 16'h7000;
    defparam add_4626_2.INIT1 = 16'h5aaa;
    defparam add_4626_2.INJECT1_0 = "NO";
    defparam add_4626_2.INJECT1_1 = "NO";
    LUT4 i49836_2_lut (.A(\buf_x[699] ), .B(\buf_x[689] ), .Z(buf_x[937])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49836_2_lut.init = 16'h6666;
    LUT4 i49850_2_lut (.A(buf_x[670]), .B(\buf_x[737] ), .Z(buf_x[938])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49850_2_lut.init = 16'h6666;
    FD1S3AX nK_b1_i9 (.D(nK_b0[8]), .CK(clock), .Q(buf_x[1002]));
    defparam nK_b1_i9.GSR = "DISABLED";
    FD1S3AX nK_b1_i8 (.D(nK_b0[7]), .CK(clock), .Q(\buf_x[727] ));
    defparam nK_b1_i8.GSR = "DISABLED";
    FD1S3AX nK_b1_i7 (.D(nK_b0[6]), .CK(clock), .Q(\buf_x[737] ));
    defparam nK_b1_i7.GSR = "DISABLED";
    FD1S3AX nK_b1_i6 (.D(nK_b0[5]), .CK(clock), .Q(\buf_x[689] ));
    defparam nK_b1_i6.GSR = "DISABLED";
    FD1S3AX nK_b1_i5 (.D(nK_b0[4]), .CK(clock), .Q(\buf_x[699] ));
    defparam nK_b1_i5.GSR = "DISABLED";
    FD1S3AX nK_b1_i4 (.D(nK_b0[3]), .CK(clock), .Q(\buf_x[651] ));
    defparam nK_b1_i4.GSR = "DISABLED";
    FD1S3AX nK_b1_i3 (.D(nK_b0[2]), .CK(clock), .Q(\buf_x[661] ));
    defparam nK_b1_i3.GSR = "DISABLED";
    FD1S3AX nK_b1_i2 (.D(nK_b0[1]), .CK(clock), .Q(\buf_x[613] ));
    defparam nK_b1_i2.GSR = "DISABLED";
    CCU2D add_2956_32 (.A0(buf_r[930]), .B0(buf_r[966]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61825), .S0(buf_x[1090]));
    defparam add_2956_32.INIT0 = 16'h5666;
    defparam add_2956_32.INIT1 = 16'h0000;
    defparam add_2956_32.INJECT1_0 = "NO";
    defparam add_2956_32.INJECT1_1 = "NO";
    CCU2D add_2956_30 (.A0(buf_r[928]), .B0(buf_r[964]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[929]), .B1(buf_r[965]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61824), .COUT(n61825), .S0(buf_x[1088]), 
          .S1(buf_x[1089]));
    defparam add_2956_30.INIT0 = 16'h5666;
    defparam add_2956_30.INIT1 = 16'h5666;
    defparam add_2956_30.INJECT1_0 = "NO";
    defparam add_2956_30.INJECT1_1 = "NO";
    CCU2D add_2956_28 (.A0(buf_r[926]), .B0(buf_r[962]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[927]), .B1(buf_r[963]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61823), .COUT(n61824), .S0(buf_x[1086]), 
          .S1(buf_x[1087]));
    defparam add_2956_28.INIT0 = 16'h5666;
    defparam add_2956_28.INIT1 = 16'h5666;
    defparam add_2956_28.INJECT1_0 = "NO";
    defparam add_2956_28.INJECT1_1 = "NO";
    CCU2D add_2956_26 (.A0(buf_r[924]), .B0(buf_r[960]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[925]), .B1(buf_r[961]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61822), .COUT(n61823), .S0(buf_x[1084]), 
          .S1(buf_x[1085]));
    defparam add_2956_26.INIT0 = 16'h5666;
    defparam add_2956_26.INIT1 = 16'h5666;
    defparam add_2956_26.INJECT1_0 = "NO";
    defparam add_2956_26.INJECT1_1 = "NO";
    CCU2D add_2956_24 (.A0(buf_r[922]), .B0(buf_r[958]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[923]), .B1(buf_r[959]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61821), .COUT(n61822), .S0(buf_x[1082]), 
          .S1(buf_x[1083]));
    defparam add_2956_24.INIT0 = 16'h5666;
    defparam add_2956_24.INIT1 = 16'h5666;
    defparam add_2956_24.INJECT1_0 = "NO";
    defparam add_2956_24.INJECT1_1 = "NO";
    CCU2D add_2956_22 (.A0(buf_r[920]), .B0(buf_r[956]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[921]), .B1(buf_r[957]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61820), .COUT(n61821), .S0(buf_x[1080]), 
          .S1(buf_x[1081]));
    defparam add_2956_22.INIT0 = 16'h5666;
    defparam add_2956_22.INIT1 = 16'h5666;
    defparam add_2956_22.INJECT1_0 = "NO";
    defparam add_2956_22.INJECT1_1 = "NO";
    CCU2D add_2956_20 (.A0(buf_r[918]), .B0(buf_r[954]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[919]), .B1(buf_r[955]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61819), .COUT(n61820), .S0(buf_x[1078]), 
          .S1(buf_x[1079]));
    defparam add_2956_20.INIT0 = 16'h5666;
    defparam add_2956_20.INIT1 = 16'h5666;
    defparam add_2956_20.INJECT1_0 = "NO";
    defparam add_2956_20.INJECT1_1 = "NO";
    CCU2D add_2956_18 (.A0(buf_r[916]), .B0(buf_r[952]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[917]), .B1(buf_r[953]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61818), .COUT(n61819), .S0(buf_x[1076]), 
          .S1(buf_x[1077]));
    defparam add_2956_18.INIT0 = 16'h5666;
    defparam add_2956_18.INIT1 = 16'h5666;
    defparam add_2956_18.INJECT1_0 = "NO";
    defparam add_2956_18.INJECT1_1 = "NO";
    CCU2D add_2956_16 (.A0(buf_r[914]), .B0(buf_r[950]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[915]), .B1(buf_r[951]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61817), .COUT(n61818), .S0(buf_x[1074]), 
          .S1(buf_x[1075]));
    defparam add_2956_16.INIT0 = 16'h5666;
    defparam add_2956_16.INIT1 = 16'h5666;
    defparam add_2956_16.INJECT1_0 = "NO";
    defparam add_2956_16.INJECT1_1 = "NO";
    CCU2D add_2956_14 (.A0(buf_r[912]), .B0(buf_r[949]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[913]), .B1(buf_r[949]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61816), .COUT(n61817), .S0(buf_x[1072]), 
          .S1(buf_x[1073]));
    defparam add_2956_14.INIT0 = 16'h5666;
    defparam add_2956_14.INIT1 = 16'h5666;
    defparam add_2956_14.INJECT1_0 = "NO";
    defparam add_2956_14.INJECT1_1 = "NO";
    CCU2D add_2956_12 (.A0(buf_r[910]), .B0(buf_r[946]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[911]), .B1(buf_r[947]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61815), .COUT(n61816), .S0(buf_x[1070]), 
          .S1(buf_x[1071]));
    defparam add_2956_12.INIT0 = 16'h5666;
    defparam add_2956_12.INIT1 = 16'h5666;
    defparam add_2956_12.INJECT1_0 = "NO";
    defparam add_2956_12.INJECT1_1 = "NO";
    CCU2D add_2956_10 (.A0(buf_r[909]), .B0(buf_r[944]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[909]), .B1(buf_r[945]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61814), .COUT(n61815), .S0(buf_x[1068]), 
          .S1(buf_x[1069]));
    defparam add_2956_10.INIT0 = 16'h5666;
    defparam add_2956_10.INIT1 = 16'h5666;
    defparam add_2956_10.INJECT1_0 = "NO";
    defparam add_2956_10.INJECT1_1 = "NO";
    CCU2D add_2956_8 (.A0(buf_r[906]), .B0(buf_r[942]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[907]), .B1(buf_r[943]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61813), .COUT(n61814), .S0(buf_x[1066]), 
          .S1(buf_x[1067]));
    defparam add_2956_8.INIT0 = 16'h5666;
    defparam add_2956_8.INIT1 = 16'h5666;
    defparam add_2956_8.INJECT1_0 = "NO";
    defparam add_2956_8.INJECT1_1 = "NO";
    CCU2D add_2956_6 (.A0(buf_r[904]), .B0(buf_r[940]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[905]), .B1(buf_r[941]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61812), .COUT(n61813), .S0(buf_x[1064]), 
          .S1(buf_x[1065]));
    defparam add_2956_6.INIT0 = 16'h5666;
    defparam add_2956_6.INIT1 = 16'h5666;
    defparam add_2956_6.INJECT1_0 = "NO";
    defparam add_2956_6.INJECT1_1 = "NO";
    CCU2D add_2956_4 (.A0(buf_r[902]), .B0(buf_r[938]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[903]), .B1(buf_r[939]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61811), .COUT(n61812), .S1(\nKLog2_c0[7] ));
    defparam add_2956_4.INIT0 = 16'h5666;
    defparam add_2956_4.INIT1 = 16'h5666;
    defparam add_2956_4.INJECT1_0 = "NO";
    defparam add_2956_4.INJECT1_1 = "NO";
    CCU2D add_2956_2 (.A0(buf_r[900]), .B0(\buf_r[936] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[901]), .B1(buf_r[937]), .C1(GND_net), 
          .D1(GND_net), .COUT(n61811));
    defparam add_2956_2.INIT0 = 16'h7000;
    defparam add_2956_2.INIT1 = 16'h5666;
    defparam add_2956_2.INJECT1_0 = "NO";
    defparam add_2956_2.INJECT1_1 = "NO";
    CCU2D add_2955_28 (.A0(buf_x[697]), .B0(buf_x[733]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[734]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61809), .S0(buf_x[965]), .S1(buf_x[966]));
    defparam add_2955_28.INIT0 = 16'h5666;
    defparam add_2955_28.INIT1 = 16'hfaaa;
    defparam add_2955_28.INJECT1_0 = "NO";
    defparam add_2955_28.INJECT1_1 = "NO";
    CCU2D add_2955_26 (.A0(buf_x[695]), .B0(buf_x[731]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[696]), .B1(buf_x[732]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61808), .COUT(n61809), .S0(buf_x[963]), 
          .S1(buf_x[964]));
    defparam add_2955_26.INIT0 = 16'h5666;
    defparam add_2955_26.INIT1 = 16'h5666;
    defparam add_2955_26.INJECT1_0 = "NO";
    defparam add_2955_26.INJECT1_1 = "NO";
    CCU2D add_2955_24 (.A0(buf_x[693]), .B0(\buf_x[737] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[694]), .B1(buf_x[730]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61807), .COUT(n61808), .S0(buf_x[961]), 
          .S1(buf_x[962]));
    defparam add_2955_24.INIT0 = 16'h5666;
    defparam add_2955_24.INIT1 = 16'h5666;
    defparam add_2955_24.INJECT1_0 = "NO";
    defparam add_2955_24.INJECT1_1 = "NO";
    CCU2D add_2955_22 (.A0(\buf_x[699] ), .B0(\buf_x[727] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[692]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61806), .COUT(n61807), .S0(buf_x[959]), 
          .S1(buf_x[960]));
    defparam add_2955_22.INIT0 = 16'h5666;
    defparam add_2955_22.INIT1 = 16'h5aaa;
    defparam add_2955_22.INJECT1_0 = "NO";
    defparam add_2955_22.INJECT1_1 = "NO";
    CCU2D add_2955_20 (.A0(\buf_x[689] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[737] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61805), .COUT(n61806), .S0(buf_x[957]), 
          .S1(buf_x[958]));
    defparam add_2955_20.INIT0 = 16'h5aaa;
    defparam add_2955_20.INIT1 = 16'hfaaa;
    defparam add_2955_20.INJECT1_0 = "NO";
    defparam add_2955_20.INJECT1_1 = "NO";
    CCU2D add_2955_18 (.A0(buf_x[723]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[699] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61804), .COUT(n61805), .S0(buf_x[955]), .S1(buf_x[956]));
    defparam add_2955_18.INIT0 = 16'hfaaa;
    defparam add_2955_18.INIT1 = 16'h5aaa;
    defparam add_2955_18.INJECT1_0 = "NO";
    defparam add_2955_18.INJECT1_1 = "NO";
    CCU2D add_2955_16 (.A0(buf_x[685]), .B0(buf_x[721]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[722]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61803), .COUT(n61804), .S0(buf_x[953]), 
          .S1(buf_x[954]));
    defparam add_2955_16.INIT0 = 16'h5666;
    defparam add_2955_16.INIT1 = 16'hfaaa;
    defparam add_2955_16.INJECT1_0 = "NO";
    defparam add_2955_16.INJECT1_1 = "NO";
    CCU2D add_2955_14 (.A0(buf_x[683]), .B0(buf_x[715]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[684]), .B1(buf_x[720]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61802), .COUT(n61803), .S0(buf_x[951]), 
          .S1(buf_x[952]));
    defparam add_2955_14.INIT0 = 16'h5666;
    defparam add_2955_14.INIT1 = 16'h5666;
    defparam add_2955_14.INJECT1_0 = "NO";
    defparam add_2955_14.INJECT1_1 = "NO";
    CCU2D add_2955_12 (.A0(buf_x[677]), .B0(buf_x[715]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[682]), .B1(buf_x[715]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61801), .COUT(n61802), .S0(buf_x[948]), 
          .S1(buf_x[950]));
    defparam add_2955_12.INIT0 = 16'h5666;
    defparam add_2955_12.INIT1 = 16'h5666;
    defparam add_2955_12.INJECT1_0 = "NO";
    defparam add_2955_12.INJECT1_1 = "NO";
    CCU2D add_2955_10 (.A0(buf_x[677]), .B0(buf_x[714]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[677]), .B1(buf_x[715]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61800), .COUT(n61801), .S0(buf_x[946]), 
          .S1(buf_x[947]));
    defparam add_2955_10.INIT0 = 16'h5666;
    defparam add_2955_10.INIT1 = 16'h5666;
    defparam add_2955_10.INJECT1_0 = "NO";
    defparam add_2955_10.INJECT1_1 = "NO";
    CCU2D add_2955_8 (.A0(buf_x[676]), .B0(buf_x[712]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[677]), .B1(buf_x[713]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61799), .COUT(n61800), .S0(buf_x[944]), 
          .S1(buf_x[945]));
    defparam add_2955_8.INIT0 = 16'h5666;
    defparam add_2955_8.INIT1 = 16'h5666;
    defparam add_2955_8.INJECT1_0 = "NO";
    defparam add_2955_8.INJECT1_1 = "NO";
    CCU2D add_2955_6 (.A0(buf_x[674]), .B0(buf_x[708]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[675]), .B1(buf_x[708]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61798), .COUT(n61799), .S0(buf_x[942]), 
          .S1(buf_x[943]));
    defparam add_2955_6.INIT0 = 16'h5666;
    defparam add_2955_6.INIT1 = 16'h5666;
    defparam add_2955_6.INJECT1_0 = "NO";
    defparam add_2955_6.INJECT1_1 = "NO";
    CCU2D add_2955_4 (.A0(buf_x[670]), .B0(buf_x[708]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[670]), .B1(buf_x[708]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61797), .COUT(n61798), .S0(buf_x[940]), 
          .S1(buf_x[941]));
    defparam add_2955_4.INIT0 = 16'h5666;
    defparam add_2955_4.INIT1 = 16'h5666;
    defparam add_2955_4.INJECT1_0 = "NO";
    defparam add_2955_4.INJECT1_1 = "NO";
    CCU2D add_2955_2 (.A0(buf_x[670]), .B0(\buf_x[737] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[737] ), .B1(\buf_x[727] ), .C1(buf_x[670]), 
          .D1(GND_net), .COUT(n61797), .S1(buf_x[939]));
    defparam add_2955_2.INIT0 = 16'h7000;
    defparam add_2955_2.INIT1 = 16'h9696;
    defparam add_2955_2.INJECT1_0 = "NO";
    defparam add_2955_2.INJECT1_1 = "NO";
    CCU2D add_2954_32 (.A0(buf_x[625]), .B0(\buf_x[661] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[626]), .B1(buf_x[662]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61794), .S0(buf_x[929]), .S1(buf_x[930]));
    defparam add_2954_32.INIT0 = 16'h5666;
    defparam add_2954_32.INIT1 = 16'h5666;
    defparam add_2954_32.INJECT1_0 = "NO";
    defparam add_2954_32.INJECT1_1 = "NO";
    CCU2D add_2954_30 (.A0(\buf_x[623] ), .B0(buf_x[659]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[624]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61793), .COUT(n61794), .S0(buf_x[927]), 
          .S1(buf_x[928]));
    defparam add_2954_30.INIT0 = 16'h5666;
    defparam add_2954_30.INIT1 = 16'h5aaa;
    defparam add_2954_30.INJECT1_0 = "NO";
    defparam add_2954_30.INJECT1_1 = "NO";
    CCU2D add_2954_28 (.A0(buf_x[621]), .B0(buf_x[657]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[658]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61792), .COUT(n61793), .S0(buf_x[925]), 
          .S1(buf_x[926]));
    defparam add_2954_28.INIT0 = 16'h5666;
    defparam add_2954_28.INIT1 = 16'hfaaa;
    defparam add_2954_28.INJECT1_0 = "NO";
    defparam add_2954_28.INJECT1_1 = "NO";
    CCU2D add_2954_26 (.A0(buf_x[619]), .B0(buf_x[655]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[620]), .B1(buf_x[656]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61791), .COUT(n61792), .S0(buf_x[923]), 
          .S1(buf_x[924]));
    defparam add_2954_26.INIT0 = 16'h5666;
    defparam add_2954_26.INIT1 = 16'h5666;
    defparam add_2954_26.INJECT1_0 = "NO";
    defparam add_2954_26.INJECT1_1 = "NO";
    CCU2D add_2954_24 (.A0(buf_x[617]), .B0(\buf_x[661] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[618]), .B1(buf_x[654]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61790), .COUT(n61791), .S0(buf_x[921]), 
          .S1(buf_x[922]));
    defparam add_2954_24.INIT0 = 16'h5666;
    defparam add_2954_24.INIT1 = 16'h5666;
    defparam add_2954_24.INJECT1_0 = "NO";
    defparam add_2954_24.INJECT1_1 = "NO";
    CCU2D add_2954_22 (.A0(\buf_x[623] ), .B0(\buf_x[651] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[616]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61789), .COUT(n61790), .S0(buf_x[919]), 
          .S1(buf_x[920]));
    defparam add_2954_22.INIT0 = 16'h5666;
    defparam add_2954_22.INIT1 = 16'h5aaa;
    defparam add_2954_22.INJECT1_0 = "NO";
    defparam add_2954_22.INJECT1_1 = "NO";
    CCU2D add_2954_20 (.A0(\buf_x[613] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[661] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61788), .COUT(n61789), .S0(buf_x[917]), 
          .S1(buf_x[918]));
    defparam add_2954_20.INIT0 = 16'h5aaa;
    defparam add_2954_20.INIT1 = 16'hfaaa;
    defparam add_2954_20.INJECT1_0 = "NO";
    defparam add_2954_20.INJECT1_1 = "NO";
    CCU2D add_2954_18 (.A0(buf_x[647]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[623] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61787), .COUT(n61788), .S0(buf_x[915]), .S1(buf_x[916]));
    defparam add_2954_18.INIT0 = 16'hfaaa;
    defparam add_2954_18.INIT1 = 16'h5aaa;
    defparam add_2954_18.INJECT1_0 = "NO";
    defparam add_2954_18.INJECT1_1 = "NO";
    CCU2D add_2954_16 (.A0(buf_x[609]), .B0(buf_x[645]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[646]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61786), .COUT(n61787), .S0(buf_x[913]), 
          .S1(buf_x[914]));
    defparam add_2954_16.INIT0 = 16'h5666;
    defparam add_2954_16.INIT1 = 16'hfaaa;
    defparam add_2954_16.INJECT1_0 = "NO";
    defparam add_2954_16.INJECT1_1 = "NO";
    CCU2D add_2954_14 (.A0(buf_x[607]), .B0(buf_x[639]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[608]), .B1(buf_x[644]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61785), .COUT(n61786), .S0(buf_x[911]), 
          .S1(buf_x[912]));
    defparam add_2954_14.INIT0 = 16'h5666;
    defparam add_2954_14.INIT1 = 16'h5666;
    defparam add_2954_14.INJECT1_0 = "NO";
    defparam add_2954_14.INJECT1_1 = "NO";
    CCU2D add_2954_12 (.A0(buf_x[601]), .B0(buf_x[639]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[606]), .B1(buf_x[639]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61784), .COUT(n61785), .S0(buf_x[908]), 
          .S1(buf_x[910]));
    defparam add_2954_12.INIT0 = 16'h5666;
    defparam add_2954_12.INIT1 = 16'h5666;
    defparam add_2954_12.INJECT1_0 = "NO";
    defparam add_2954_12.INJECT1_1 = "NO";
    CCU2D add_2954_10 (.A0(buf_x[601]), .B0(buf_x[638]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[601]), .B1(buf_x[639]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61783), .COUT(n61784), .S0(buf_x[906]), 
          .S1(buf_x[907]));
    defparam add_2954_10.INIT0 = 16'h5666;
    defparam add_2954_10.INIT1 = 16'h5666;
    defparam add_2954_10.INJECT1_0 = "NO";
    defparam add_2954_10.INJECT1_1 = "NO";
    CCU2D add_2954_8 (.A0(buf_x[600]), .B0(buf_x[636]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[601]), .B1(buf_x[637]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61782), .COUT(n61783), .S0(buf_x[904]), 
          .S1(buf_x[905]));
    defparam add_2954_8.INIT0 = 16'h5666;
    defparam add_2954_8.INIT1 = 16'h5666;
    defparam add_2954_8.INJECT1_0 = "NO";
    defparam add_2954_8.INJECT1_1 = "NO";
    CCU2D add_2954_6 (.A0(buf_x[598]), .B0(buf_x[632]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[599]), .B1(buf_x[632]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61781), .COUT(n61782), .S0(buf_x[902]), 
          .S1(buf_x[903]));
    defparam add_2954_6.INIT0 = 16'h5666;
    defparam add_2954_6.INIT1 = 16'h5666;
    defparam add_2954_6.INJECT1_0 = "NO";
    defparam add_2954_6.INJECT1_1 = "NO";
    CCU2D add_2954_4 (.A0(buf_x[594]), .B0(buf_x[632]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[594]), .B1(buf_x[632]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61780), .COUT(n61781), .S0(buf_x[900]), 
          .S1(buf_x[901]));
    defparam add_2954_4.INIT0 = 16'h5666;
    defparam add_2954_4.INIT1 = 16'h5666;
    defparam add_2954_4.INJECT1_0 = "NO";
    defparam add_2954_4.INJECT1_1 = "NO";
    CCU2D add_2954_2 (.A0(buf_x[594]), .B0(\buf_x[661] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[661] ), .B1(\buf_x[651] ), .C1(buf_x[594]), 
          .D1(GND_net), .COUT(n61780));
    defparam add_2954_2.INIT0 = 16'h7000;
    defparam add_2954_2.INIT1 = 16'h9696;
    defparam add_2954_2.INJECT1_0 = "NO";
    defparam add_2954_2.INJECT1_1 = "NO";
    CCU2D add_4602_20 (.A0(\buf_x[737] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[727] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61764), .S0(buf_x[733]), .S1(buf_x[734]));
    defparam add_4602_20.INIT0 = 16'h5aaa;
    defparam add_4602_20.INIT1 = 16'hfaaa;
    defparam add_4602_20.INJECT1_0 = "NO";
    defparam add_4602_20.INJECT1_1 = "NO";
    CCU2D add_4602_18 (.A0(\buf_x[737] ), .B0(\buf_x[727] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[727] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61763), .COUT(n61764), .S0(buf_x[731]), 
          .S1(buf_x[732]));
    defparam add_4602_18.INIT0 = 16'h5666;
    defparam add_4602_18.INIT1 = 16'hfaaa;
    defparam add_4602_18.INJECT1_0 = "NO";
    defparam add_4602_18.INJECT1_1 = "NO";
    CCU2D add_4602_16 (.A0(\buf_x[737] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[737] ), .B1(\buf_x[727] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61762), .COUT(n61763), .S1(buf_x[730]));
    defparam add_4602_16.INIT0 = 16'h5aaa;
    defparam add_4602_16.INIT1 = 16'h5666;
    defparam add_4602_16.INJECT1_0 = "NO";
    defparam add_4602_16.INJECT1_1 = "NO";
    CCU2D add_4602_14 (.A0(\buf_x[727] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61761), .COUT(n61762));
    defparam add_4602_14.INIT0 = 16'hfaaa;
    defparam add_4602_14.INIT1 = 16'hf000;
    defparam add_4602_14.INJECT1_0 = "NO";
    defparam add_4602_14.INJECT1_1 = "NO";
    CCU2D add_4602_12 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[737] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61760), .COUT(n61761));
    defparam add_4602_12.INIT0 = 16'hf000;
    defparam add_4602_12.INIT1 = 16'h5aaa;
    defparam add_4602_12.INJECT1_0 = "NO";
    defparam add_4602_12.INJECT1_1 = "NO";
    CCU2D add_4602_10 (.A0(\buf_x[727] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61759), .COUT(n61760), .S0(buf_x[722]), .S1(buf_x[723]));
    defparam add_4602_10.INIT0 = 16'hfaaa;
    defparam add_4602_10.INIT1 = 16'hf000;
    defparam add_4602_10.INJECT1_0 = "NO";
    defparam add_4602_10.INJECT1_1 = "NO";
    CCU2D add_4602_8 (.A0(\buf_x[727] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[737] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61758), .COUT(n61759), .S0(buf_x[720]), .S1(buf_x[721]));
    defparam add_4602_8.INIT0 = 16'hfaaa;
    defparam add_4602_8.INIT1 = 16'h5aaa;
    defparam add_4602_8.INJECT1_0 = "NO";
    defparam add_4602_8.INJECT1_1 = "NO";
    CCU2D add_4602_6 (.A0(\buf_x[737] ), .B0(\buf_x[727] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[737] ), .B1(\buf_x[727] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61757), .COUT(n61758), .S0(buf_x[714]), 
          .S1(buf_x[715]));
    defparam add_4602_6.INIT0 = 16'h5666;
    defparam add_4602_6.INIT1 = 16'h5666;
    defparam add_4602_6.INJECT1_0 = "NO";
    defparam add_4602_6.INJECT1_1 = "NO";
    CCU2D add_4602_4 (.A0(\buf_x[727] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[737] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61756), .COUT(n61757), .S0(buf_x[712]), .S1(buf_x[713]));
    defparam add_4602_4.INIT0 = 16'hfaaa;
    defparam add_4602_4.INIT1 = 16'h5aaa;
    defparam add_4602_4.INJECT1_0 = "NO";
    defparam add_4602_4.INJECT1_1 = "NO";
    CCU2D add_4602_2 (.A0(\buf_x[737] ), .B0(\buf_x[727] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[737] ), .B1(\buf_x[727] ), .C1(GND_net), 
          .D1(GND_net), .COUT(n61756), .S1(buf_x[708]));
    defparam add_4602_2.INIT0 = 16'h7000;
    defparam add_4602_2.INIT1 = 16'h5666;
    defparam add_4602_2.INJECT1_0 = "NO";
    defparam add_4602_2.INJECT1_1 = "NO";
    CCU2D add_4600_24 (.A0(\buf_x[661] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[661] ), .B1(\buf_x[651] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61749), .S1(buf_x[662]));
    defparam add_4600_24.INIT0 = 16'h5aaa;
    defparam add_4600_24.INIT1 = 16'h5666;
    defparam add_4600_24.INJECT1_0 = "NO";
    defparam add_4600_24.INJECT1_1 = "NO";
    CCU2D add_4600_22 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61748), 
          .COUT(n61749), .S0(buf_x[659]));
    defparam add_4600_22.INIT0 = 16'hf000;
    defparam add_4600_22.INIT1 = 16'hf000;
    defparam add_4600_22.INJECT1_0 = "NO";
    defparam add_4600_22.INJECT1_1 = "NO";
    CCU2D add_4600_20 (.A0(\buf_x[661] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[651] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61747), .COUT(n61748), .S0(buf_x[657]), 
          .S1(buf_x[658]));
    defparam add_4600_20.INIT0 = 16'h5aaa;
    defparam add_4600_20.INIT1 = 16'hfaaa;
    defparam add_4600_20.INJECT1_0 = "NO";
    defparam add_4600_20.INJECT1_1 = "NO";
    CCU2D add_4600_18 (.A0(\buf_x[661] ), .B0(\buf_x[651] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[651] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61746), .COUT(n61747), .S0(buf_x[655]), 
          .S1(buf_x[656]));
    defparam add_4600_18.INIT0 = 16'h5666;
    defparam add_4600_18.INIT1 = 16'hfaaa;
    defparam add_4600_18.INJECT1_0 = "NO";
    defparam add_4600_18.INJECT1_1 = "NO";
    CCU2D add_4600_16 (.A0(\buf_x[661] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[661] ), .B1(\buf_x[651] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61745), .COUT(n61746), .S1(buf_x[654]));
    defparam add_4600_16.INIT0 = 16'h5aaa;
    defparam add_4600_16.INIT1 = 16'h5666;
    defparam add_4600_16.INJECT1_0 = "NO";
    defparam add_4600_16.INJECT1_1 = "NO";
    CCU2D add_4600_14 (.A0(\buf_x[651] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61744), .COUT(n61745));
    defparam add_4600_14.INIT0 = 16'hfaaa;
    defparam add_4600_14.INIT1 = 16'hf000;
    defparam add_4600_14.INJECT1_0 = "NO";
    defparam add_4600_14.INJECT1_1 = "NO";
    CCU2D add_4600_12 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[661] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61743), .COUT(n61744));
    defparam add_4600_12.INIT0 = 16'hf000;
    defparam add_4600_12.INIT1 = 16'h5aaa;
    defparam add_4600_12.INJECT1_0 = "NO";
    defparam add_4600_12.INJECT1_1 = "NO";
    CCU2D add_4600_10 (.A0(\buf_x[651] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61742), .COUT(n61743), .S0(buf_x[646]), .S1(buf_x[647]));
    defparam add_4600_10.INIT0 = 16'hfaaa;
    defparam add_4600_10.INIT1 = 16'hf000;
    defparam add_4600_10.INJECT1_0 = "NO";
    defparam add_4600_10.INJECT1_1 = "NO";
    CCU2D add_4600_8 (.A0(\buf_x[651] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[661] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61741), .COUT(n61742), .S0(buf_x[644]), .S1(buf_x[645]));
    defparam add_4600_8.INIT0 = 16'hfaaa;
    defparam add_4600_8.INIT1 = 16'h5aaa;
    defparam add_4600_8.INJECT1_0 = "NO";
    defparam add_4600_8.INJECT1_1 = "NO";
    CCU2D add_4600_6 (.A0(\buf_x[661] ), .B0(\buf_x[651] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[661] ), .B1(\buf_x[651] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61740), .COUT(n61741), .S0(buf_x[638]), 
          .S1(buf_x[639]));
    defparam add_4600_6.INIT0 = 16'h5666;
    defparam add_4600_6.INIT1 = 16'h5666;
    defparam add_4600_6.INJECT1_0 = "NO";
    defparam add_4600_6.INJECT1_1 = "NO";
    CCU2D add_4600_4 (.A0(\buf_x[651] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[661] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61739), .COUT(n61740), .S0(buf_x[636]), .S1(buf_x[637]));
    defparam add_4600_4.INIT0 = 16'hfaaa;
    defparam add_4600_4.INIT1 = 16'h5aaa;
    defparam add_4600_4.INJECT1_0 = "NO";
    defparam add_4600_4.INJECT1_1 = "NO";
    CCU2D add_4600_2 (.A0(\buf_x[661] ), .B0(\buf_x[651] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[661] ), .B1(\buf_x[651] ), .C1(GND_net), 
          .D1(GND_net), .COUT(n61739), .S1(buf_x[632]));
    defparam add_4600_2.INIT0 = 16'h7000;
    defparam add_4600_2.INIT1 = 16'h5666;
    defparam add_4600_2.INJECT1_0 = "NO";
    defparam add_4600_2.INJECT1_1 = "NO";
    LUT4 i49857_2_lut (.A(buf_x[1064]), .B(buf_x[1100]), .Z(\nKLog2_c0[8] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49857_2_lut.init = 16'h6666;
    CCU2D add_4599_26 (.A0(\buf_x[613] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[623] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61707), .S0(buf_x[625]), .S1(buf_x[626]));
    defparam add_4599_26.INIT0 = 16'hfaaa;
    defparam add_4599_26.INIT1 = 16'h5aaa;
    defparam add_4599_26.INJECT1_0 = "NO";
    defparam add_4599_26.INJECT1_1 = "NO";
    CCU2D add_4599_24 (.A0(\buf_x[623] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[623] ), .B1(\buf_x[613] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61706), .COUT(n61707), .S1(buf_x[624]));
    defparam add_4599_24.INIT0 = 16'h5aaa;
    defparam add_4599_24.INIT1 = 16'h5666;
    defparam add_4599_24.INJECT1_0 = "NO";
    defparam add_4599_24.INJECT1_1 = "NO";
    CCU2D add_4599_22 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61705), 
          .COUT(n61706), .S0(buf_x[621]));
    defparam add_4599_22.INIT0 = 16'hf000;
    defparam add_4599_22.INIT1 = 16'hf000;
    defparam add_4599_22.INJECT1_0 = "NO";
    defparam add_4599_22.INJECT1_1 = "NO";
    CCU2D add_4599_20 (.A0(\buf_x[623] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[613] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61704), .COUT(n61705), .S0(buf_x[619]), 
          .S1(buf_x[620]));
    defparam add_4599_20.INIT0 = 16'h5aaa;
    defparam add_4599_20.INIT1 = 16'hfaaa;
    defparam add_4599_20.INJECT1_0 = "NO";
    defparam add_4599_20.INJECT1_1 = "NO";
    CCU2D add_4599_18 (.A0(\buf_x[623] ), .B0(\buf_x[613] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[613] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61703), .COUT(n61704), .S0(buf_x[617]), 
          .S1(buf_x[618]));
    defparam add_4599_18.INIT0 = 16'h5666;
    defparam add_4599_18.INIT1 = 16'hfaaa;
    defparam add_4599_18.INJECT1_0 = "NO";
    defparam add_4599_18.INJECT1_1 = "NO";
    CCU2D add_4599_16 (.A0(\buf_x[623] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[623] ), .B1(\buf_x[613] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61702), .COUT(n61703), .S1(buf_x[616]));
    defparam add_4599_16.INIT0 = 16'h5aaa;
    defparam add_4599_16.INIT1 = 16'h5666;
    defparam add_4599_16.INJECT1_0 = "NO";
    defparam add_4599_16.INJECT1_1 = "NO";
    CCU2D add_4599_14 (.A0(\buf_x[613] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61701), .COUT(n61702));
    defparam add_4599_14.INIT0 = 16'hfaaa;
    defparam add_4599_14.INIT1 = 16'hf000;
    defparam add_4599_14.INJECT1_0 = "NO";
    defparam add_4599_14.INJECT1_1 = "NO";
    CCU2D add_4599_12 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[623] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61700), .COUT(n61701));
    defparam add_4599_12.INIT0 = 16'hf000;
    defparam add_4599_12.INIT1 = 16'h5aaa;
    defparam add_4599_12.INJECT1_0 = "NO";
    defparam add_4599_12.INJECT1_1 = "NO";
    CCU2D add_4599_10 (.A0(\buf_x[613] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61699), .COUT(n61700), .S0(buf_x[608]), .S1(buf_x[609]));
    defparam add_4599_10.INIT0 = 16'hfaaa;
    defparam add_4599_10.INIT1 = 16'hf000;
    defparam add_4599_10.INJECT1_0 = "NO";
    defparam add_4599_10.INJECT1_1 = "NO";
    CCU2D add_4599_8 (.A0(\buf_x[613] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[623] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61698), .COUT(n61699), .S0(buf_x[606]), .S1(buf_x[607]));
    defparam add_4599_8.INIT0 = 16'hfaaa;
    defparam add_4599_8.INIT1 = 16'h5aaa;
    defparam add_4599_8.INJECT1_0 = "NO";
    defparam add_4599_8.INJECT1_1 = "NO";
    CCU2D add_4599_6 (.A0(\buf_x[623] ), .B0(\buf_x[613] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[623] ), .B1(\buf_x[613] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61697), .COUT(n61698), .S0(buf_x[600]), 
          .S1(buf_x[601]));
    defparam add_4599_6.INIT0 = 16'h5666;
    defparam add_4599_6.INIT1 = 16'h5666;
    defparam add_4599_6.INJECT1_0 = "NO";
    defparam add_4599_6.INJECT1_1 = "NO";
    CCU2D add_4599_4 (.A0(\buf_x[613] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[623] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61696), .COUT(n61697), .S0(buf_x[598]), .S1(buf_x[599]));
    defparam add_4599_4.INIT0 = 16'hfaaa;
    defparam add_4599_4.INIT1 = 16'h5aaa;
    defparam add_4599_4.INJECT1_0 = "NO";
    defparam add_4599_4.INJECT1_1 = "NO";
    CCU2D add_4599_2 (.A0(\buf_x[623] ), .B0(\buf_x[613] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[623] ), .B1(\buf_x[613] ), .C1(GND_net), 
          .D1(GND_net), .COUT(n61696), .S1(buf_x[594]));
    defparam add_4599_2.INIT0 = 16'h7000;
    defparam add_4599_2.INIT1 = 16'h5666;
    defparam add_4599_2.INJECT1_0 = "NO";
    defparam add_4599_2.INJECT1_1 = "NO";
    CCU2D add_4696_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61498), 
          .S0(buf_x[697]));
    defparam add_4696_cout.INIT0 = 16'h0000;
    defparam add_4696_cout.INIT1 = 16'h0000;
    defparam add_4696_cout.INJECT1_0 = "NO";
    defparam add_4696_cout.INJECT1_1 = "NO";
    CCU2D add_4696_20 (.A0(\buf_x[699] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[689] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61497), .COUT(n61498), .S0(buf_x[695]), 
          .S1(buf_x[696]));
    defparam add_4696_20.INIT0 = 16'h5aaa;
    defparam add_4696_20.INIT1 = 16'hfaaa;
    defparam add_4696_20.INJECT1_0 = "NO";
    defparam add_4696_20.INJECT1_1 = "NO";
    CCU2D add_4696_18 (.A0(\buf_x[699] ), .B0(\buf_x[689] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[689] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61496), .COUT(n61497), .S0(buf_x[693]), 
          .S1(buf_x[694]));
    defparam add_4696_18.INIT0 = 16'h5666;
    defparam add_4696_18.INIT1 = 16'hfaaa;
    defparam add_4696_18.INJECT1_0 = "NO";
    defparam add_4696_18.INJECT1_1 = "NO";
    CCU2D add_4696_16 (.A0(\buf_x[699] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[699] ), .B1(\buf_x[689] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61495), .COUT(n61496), .S1(buf_x[692]));
    defparam add_4696_16.INIT0 = 16'h5aaa;
    defparam add_4696_16.INIT1 = 16'h5666;
    defparam add_4696_16.INJECT1_0 = "NO";
    defparam add_4696_16.INJECT1_1 = "NO";
    CCU2D add_4696_14 (.A0(\buf_x[689] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61494), .COUT(n61495));
    defparam add_4696_14.INIT0 = 16'hfaaa;
    defparam add_4696_14.INIT1 = 16'hf000;
    defparam add_4696_14.INJECT1_0 = "NO";
    defparam add_4696_14.INJECT1_1 = "NO";
    CCU2D add_4696_12 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[699] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61493), .COUT(n61494));
    defparam add_4696_12.INIT0 = 16'hf000;
    defparam add_4696_12.INIT1 = 16'h5aaa;
    defparam add_4696_12.INJECT1_0 = "NO";
    defparam add_4696_12.INJECT1_1 = "NO";
    CCU2D add_4696_10 (.A0(\buf_x[689] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61492), .COUT(n61493), .S0(buf_x[684]), .S1(buf_x[685]));
    defparam add_4696_10.INIT0 = 16'hfaaa;
    defparam add_4696_10.INIT1 = 16'hf000;
    defparam add_4696_10.INJECT1_0 = "NO";
    defparam add_4696_10.INJECT1_1 = "NO";
    CCU2D add_4696_8 (.A0(\buf_x[689] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[699] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61491), .COUT(n61492), .S0(buf_x[682]), .S1(buf_x[683]));
    defparam add_4696_8.INIT0 = 16'hfaaa;
    defparam add_4696_8.INIT1 = 16'h5aaa;
    defparam add_4696_8.INJECT1_0 = "NO";
    defparam add_4696_8.INJECT1_1 = "NO";
    CCU2D add_4696_6 (.A0(\buf_x[699] ), .B0(\buf_x[689] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[699] ), .B1(\buf_x[689] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61490), .COUT(n61491), .S0(buf_x[676]), 
          .S1(buf_x[677]));
    defparam add_4696_6.INIT0 = 16'h5666;
    defparam add_4696_6.INIT1 = 16'h5666;
    defparam add_4696_6.INJECT1_0 = "NO";
    defparam add_4696_6.INJECT1_1 = "NO";
    CCU2D add_4696_4 (.A0(\buf_x[689] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\buf_x[699] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61489), .COUT(n61490), .S0(buf_x[674]), .S1(buf_x[675]));
    defparam add_4696_4.INIT0 = 16'hfaaa;
    defparam add_4696_4.INIT1 = 16'h5aaa;
    defparam add_4696_4.INJECT1_0 = "NO";
    defparam add_4696_4.INJECT1_1 = "NO";
    CCU2D add_4696_2 (.A0(\buf_x[699] ), .B0(\buf_x[689] ), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_x[699] ), .B1(\buf_x[689] ), .C1(GND_net), 
          .D1(GND_net), .COUT(n61489), .S1(buf_x[670]));
    defparam add_4696_2.INIT0 = 16'h7000;
    defparam add_4696_2.INIT1 = 16'h5666;
    defparam add_4696_2.INJECT1_0 = "NO";
    defparam add_4696_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \mult_clk(12,10,true,false,0,3) 
//

module \mult_clk(12,10,true,false,0,3)  (\nX_a1[0] , clock, \eX_x[11] , 
            \buf_x[463] , \buf_x[437] , \buf_x[436] , \buf_x[435] , 
            \buf_x[434] , \nX_a0[35] , \nX_a0[34] , \nX_a0[33] , \nX_a0[32] , 
            \nX_a0[31] , \nX_a0[30] , \nX_a0[29] , \nX_a0[28] , \nX_a0[27] , 
            \nX_a0[26] , \nX_a0[25] , \nX_a0[24] , \nX_a1[23] , \nX_a0[23] , 
            \nX_a1[22] , \nX_a0[22] , \nX_a1[21] , \nX_a0[21] , \nX_a1[20] , 
            \nX_a0[20] , \nX_a1[19] , \nX_a0[19] , \nX_a1[18] , \nX_a0[18] , 
            \nX_a1[17] , \nX_a0[17] , \nX_a1[16] , \nX_a0[16] , \nX_a1[15] , 
            \nX_a0[15] , \nX_a1[14] , \nX_a0[14] , \nX_a1[13] , \nX_a0[13] , 
            \nX_a1[12] , \nX_a0[12] , \nX_a1[11] , \nX_a0[11] , \nX_a1[10] , 
            \nX_a0[10] , \nX_a1[9] , \nX_a0[9] , \nX_a1[8] , \buf_x[471] , 
            \nX_a1[7] , \buf_x[470] , \nX_a1[6] , \buf_x[469] , \nX_a1[5] , 
            \buf_x[468] , \nX_a1[4] , \buf_x[467] , \nX_a1[3] , \buf_x[466] , 
            \nX_a1[2] , \buf_x[465] , \nX_a1[1] , \buf_x[464] , GND_net, 
            \nK0_b0[21] , \nK0_b0[19] , \nK0_b0[20] , \nK0_b0[17] , 
            \nK0_b0[18] , \nK0_b0[15] , \nK0_b0[16] , \nK0_b0[13] , 
            \nK0_b0[14] , \nK0_b0[12] );
    output \nX_a1[0] ;
    input clock;
    input \eX_x[11] ;
    input \buf_x[463] ;
    output \buf_x[437] ;
    output \buf_x[436] ;
    output \buf_x[435] ;
    output \buf_x[434] ;
    input \nX_a0[35] ;
    input \nX_a0[34] ;
    input \nX_a0[33] ;
    input \nX_a0[32] ;
    input \nX_a0[31] ;
    input \nX_a0[30] ;
    input \nX_a0[29] ;
    input \nX_a0[28] ;
    input \nX_a0[27] ;
    input \nX_a0[26] ;
    input \nX_a0[25] ;
    input \nX_a0[24] ;
    output \nX_a1[23] ;
    input \nX_a0[23] ;
    output \nX_a1[22] ;
    input \nX_a0[22] ;
    output \nX_a1[21] ;
    input \nX_a0[21] ;
    output \nX_a1[20] ;
    input \nX_a0[20] ;
    output \nX_a1[19] ;
    input \nX_a0[19] ;
    output \nX_a1[18] ;
    input \nX_a0[18] ;
    output \nX_a1[17] ;
    input \nX_a0[17] ;
    output \nX_a1[16] ;
    input \nX_a0[16] ;
    output \nX_a1[15] ;
    input \nX_a0[15] ;
    output \nX_a1[14] ;
    input \nX_a0[14] ;
    output \nX_a1[13] ;
    input \nX_a0[13] ;
    output \nX_a1[12] ;
    input \nX_a0[12] ;
    output \nX_a1[11] ;
    input \nX_a0[11] ;
    output \nX_a1[10] ;
    input \nX_a0[10] ;
    output \nX_a1[9] ;
    input \nX_a0[9] ;
    output \nX_a1[8] ;
    input \buf_x[471] ;
    output \nX_a1[7] ;
    input \buf_x[470] ;
    output \nX_a1[6] ;
    input \buf_x[469] ;
    output \nX_a1[5] ;
    input \buf_x[468] ;
    output \nX_a1[4] ;
    input \buf_x[467] ;
    output \nX_a1[3] ;
    input \buf_x[466] ;
    output \nX_a1[2] ;
    input \buf_x[465] ;
    output \nX_a1[1] ;
    input \buf_x[464] ;
    input GND_net;
    output \nK0_b0[21] ;
    output \nK0_b0[19] ;
    output \nK0_b0[20] ;
    output \nK0_b0[17] ;
    output \nK0_b0[18] ;
    output \nK0_b0[15] ;
    output \nK0_b0[16] ;
    output \nK0_b0[13] ;
    output \nK0_b0[14] ;
    output \nK0_b0[12] ;
    
    wire [482:0]buf_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [482:0]buf_r;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(337[10:15])
    
    wire n61737, n61736, n61735, n61734, n61733, n61732, n61731, 
        n61730, n61729, n61728, n61727, n61726, n61725, n61722, 
        n61721, n61720, n61719, n61718, n61717, n61716, n61715, 
        n61714, n61713, n61712, n61711, n61710;
    
    FD1S3IX nX_a1_i0 (.D(\buf_x[463] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[0] ));
    defparam nX_a1_i0.GSR = "DISABLED";
    FD1S3AX buf_r_391__77 (.D(buf_x[268]), .CK(clock), .Q(buf_x[446]));
    defparam buf_r_391__77.GSR = "DISABLED";
    FD1S3AX buf_r_389__79 (.D(buf_x[389]), .CK(clock), .Q(buf_x[444]));
    defparam buf_r_389__79.GSR = "DISABLED";
    FD1S3AX buf_r_388__80 (.D(buf_x[388]), .CK(clock), .Q(buf_x[443]));
    defparam buf_r_388__80.GSR = "DISABLED";
    FD1S3AX buf_r_387__81 (.D(buf_x[387]), .CK(clock), .Q(buf_x[442]));
    defparam buf_r_387__81.GSR = "DISABLED";
    FD1S3AX buf_r_386__82 (.D(buf_x[386]), .CK(clock), .Q(buf_x[441]));
    defparam buf_r_386__82.GSR = "DISABLED";
    FD1S3AX buf_r_385__83 (.D(buf_x[385]), .CK(clock), .Q(buf_x[440]));
    defparam buf_r_385__83.GSR = "DISABLED";
    FD1S3AX buf_r_384__84 (.D(buf_x[384]), .CK(clock), .Q(buf_x[439]));
    defparam buf_r_384__84.GSR = "DISABLED";
    FD1S3AX buf_r_383__85 (.D(buf_x[383]), .CK(clock), .Q(buf_x[438]));
    defparam buf_r_383__85.GSR = "DISABLED";
    FD1S3AX buf_r_382__86 (.D(buf_x[382]), .CK(clock), .Q(\buf_x[437] ));
    defparam buf_r_382__86.GSR = "DISABLED";
    FD1S3AX buf_r_381__87 (.D(buf_x[381]), .CK(clock), .Q(\buf_x[436] ));
    defparam buf_r_381__87.GSR = "DISABLED";
    FD1S3AX buf_r_380__88 (.D(buf_x[380]), .CK(clock), .Q(\buf_x[435] ));
    defparam buf_r_380__88.GSR = "DISABLED";
    FD1S3AX buf_r_379__89 (.D(buf_x[379]), .CK(clock), .Q(\buf_x[434] ));
    defparam buf_r_379__89.GSR = "DISABLED";
    FD1S3AX buf_r_377__91 (.D(buf_x[377]), .CK(clock), .Q(buf_r[377]));
    defparam buf_r_377__91.GSR = "DISABLED";
    FD1S3AX buf_r_376__92 (.D(buf_x[376]), .CK(clock), .Q(buf_r[376]));
    defparam buf_r_376__92.GSR = "DISABLED";
    FD1S3AX buf_r_375__93 (.D(buf_x[375]), .CK(clock), .Q(buf_r[375]));
    defparam buf_r_375__93.GSR = "DISABLED";
    FD1S3AX buf_r_374__94 (.D(buf_x[374]), .CK(clock), .Q(buf_r[374]));
    defparam buf_r_374__94.GSR = "DISABLED";
    FD1S3AX buf_r_373__95 (.D(buf_x[373]), .CK(clock), .Q(buf_r[373]));
    defparam buf_r_373__95.GSR = "DISABLED";
    FD1S3AX buf_r_372__96 (.D(buf_x[372]), .CK(clock), .Q(buf_r[372]));
    defparam buf_r_372__96.GSR = "DISABLED";
    FD1S3AX buf_r_371__97 (.D(buf_x[371]), .CK(clock), .Q(buf_r[371]));
    defparam buf_r_371__97.GSR = "DISABLED";
    FD1S3AX buf_r_370__98 (.D(buf_x[370]), .CK(clock), .Q(buf_r[370]));
    defparam buf_r_370__98.GSR = "DISABLED";
    FD1S3AX buf_r_369__99 (.D(buf_x[369]), .CK(clock), .Q(buf_r[369]));
    defparam buf_r_369__99.GSR = "DISABLED";
    FD1S3AX buf_r_368__100 (.D(buf_x[368]), .CK(clock), .Q(buf_r[368]));
    defparam buf_r_368__100.GSR = "DISABLED";
    FD1S3AX buf_r_367__101 (.D(buf_x[367]), .CK(clock), .Q(buf_r[367]));
    defparam buf_r_367__101.GSR = "DISABLED";
    FD1S3AX buf_r_366__102 (.D(buf_x[366]), .CK(clock), .Q(buf_r[366]));
    defparam buf_r_366__102.GSR = "DISABLED";
    FD1S3AX buf_r_365__103 (.D(buf_x[365]), .CK(clock), .Q(buf_r[365]));
    defparam buf_r_365__103.GSR = "DISABLED";
    FD1S3AX buf_r_364__104 (.D(buf_x[364]), .CK(clock), .Q(buf_r[364]));
    defparam buf_r_364__104.GSR = "DISABLED";
    FD1S3AX buf_r_363__105 (.D(buf_x[363]), .CK(clock), .Q(buf_r[363]));
    defparam buf_r_363__105.GSR = "DISABLED";
    FD1S3AX buf_r_357__111 (.D(buf_x[357]), .CK(clock), .Q(buf_r[357]));
    defparam buf_r_357__111.GSR = "DISABLED";
    FD1S3AX buf_r_356__112 (.D(buf_x[356]), .CK(clock), .Q(buf_r[356]));
    defparam buf_r_356__112.GSR = "DISABLED";
    FD1S3AX buf_r_355__113 (.D(buf_x[355]), .CK(clock), .Q(buf_r[355]));
    defparam buf_r_355__113.GSR = "DISABLED";
    FD1S3AX buf_r_354__114 (.D(buf_x[354]), .CK(clock), .Q(buf_r[354]));
    defparam buf_r_354__114.GSR = "DISABLED";
    FD1S3AX buf_r_353__115 (.D(buf_x[353]), .CK(clock), .Q(buf_r[353]));
    defparam buf_r_353__115.GSR = "DISABLED";
    FD1S3AX buf_r_352__116 (.D(buf_x[352]), .CK(clock), .Q(buf_r[352]));
    defparam buf_r_352__116.GSR = "DISABLED";
    FD1S3AX buf_r_351__117 (.D(buf_x[351]), .CK(clock), .Q(buf_r[351]));
    defparam buf_r_351__117.GSR = "DISABLED";
    FD1S3AX buf_r_350__118 (.D(buf_x[350]), .CK(clock), .Q(buf_r[350]));
    defparam buf_r_350__118.GSR = "DISABLED";
    FD1S3AX buf_r_349__119 (.D(buf_x[349]), .CK(clock), .Q(buf_r[349]));
    defparam buf_r_349__119.GSR = "DISABLED";
    LUT4 i49847_2_lut (.A(buf_x[380]), .B(buf_x[379]), .Z(buf_x[363])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49847_2_lut.init = 16'h6666;
    FD1S3AX nX_a1_i35 (.D(\nX_a0[35] ), .CK(clock), .Q(buf_x[268]));
    defparam nX_a1_i35.GSR = "DISABLED";
    FD1S3AX nX_a1_i34 (.D(\nX_a0[34] ), .CK(clock), .Q(buf_x[389]));
    defparam nX_a1_i34.GSR = "DISABLED";
    FD1S3AX nX_a1_i33 (.D(\nX_a0[33] ), .CK(clock), .Q(buf_x[388]));
    defparam nX_a1_i33.GSR = "DISABLED";
    FD1S3AX nX_a1_i32 (.D(\nX_a0[32] ), .CK(clock), .Q(buf_x[387]));
    defparam nX_a1_i32.GSR = "DISABLED";
    FD1S3AX nX_a1_i31 (.D(\nX_a0[31] ), .CK(clock), .Q(buf_x[386]));
    defparam nX_a1_i31.GSR = "DISABLED";
    FD1S3AX nX_a1_i30 (.D(\nX_a0[30] ), .CK(clock), .Q(buf_x[385]));
    defparam nX_a1_i30.GSR = "DISABLED";
    FD1S3AX nX_a1_i29 (.D(\nX_a0[29] ), .CK(clock), .Q(buf_x[384]));
    defparam nX_a1_i29.GSR = "DISABLED";
    FD1S3AX nX_a1_i28 (.D(\nX_a0[28] ), .CK(clock), .Q(buf_x[383]));
    defparam nX_a1_i28.GSR = "DISABLED";
    FD1S3AX nX_a1_i27 (.D(\nX_a0[27] ), .CK(clock), .Q(buf_x[382]));
    defparam nX_a1_i27.GSR = "DISABLED";
    FD1S3AX nX_a1_i26 (.D(\nX_a0[26] ), .CK(clock), .Q(buf_x[381]));
    defparam nX_a1_i26.GSR = "DISABLED";
    FD1S3AX nX_a1_i25 (.D(\nX_a0[25] ), .CK(clock), .Q(buf_x[380]));
    defparam nX_a1_i25.GSR = "DISABLED";
    FD1S3AX nX_a1_i24 (.D(\nX_a0[24] ), .CK(clock), .Q(buf_x[379]));
    defparam nX_a1_i24.GSR = "DISABLED";
    FD1S3AX nX_a1_i23 (.D(\nX_a0[23] ), .CK(clock), .Q(\nX_a1[23] ));
    defparam nX_a1_i23.GSR = "DISABLED";
    FD1S3AX nX_a1_i22 (.D(\nX_a0[22] ), .CK(clock), .Q(\nX_a1[22] ));
    defparam nX_a1_i22.GSR = "DISABLED";
    FD1S3AX nX_a1_i21 (.D(\nX_a0[21] ), .CK(clock), .Q(\nX_a1[21] ));
    defparam nX_a1_i21.GSR = "DISABLED";
    FD1S3AX nX_a1_i20 (.D(\nX_a0[20] ), .CK(clock), .Q(\nX_a1[20] ));
    defparam nX_a1_i20.GSR = "DISABLED";
    FD1S3AX nX_a1_i19 (.D(\nX_a0[19] ), .CK(clock), .Q(\nX_a1[19] ));
    defparam nX_a1_i19.GSR = "DISABLED";
    FD1S3AX nX_a1_i18 (.D(\nX_a0[18] ), .CK(clock), .Q(\nX_a1[18] ));
    defparam nX_a1_i18.GSR = "DISABLED";
    FD1S3AX nX_a1_i17 (.D(\nX_a0[17] ), .CK(clock), .Q(\nX_a1[17] ));
    defparam nX_a1_i17.GSR = "DISABLED";
    FD1S3AX nX_a1_i16 (.D(\nX_a0[16] ), .CK(clock), .Q(\nX_a1[16] ));
    defparam nX_a1_i16.GSR = "DISABLED";
    FD1S3AX nX_a1_i15 (.D(\nX_a0[15] ), .CK(clock), .Q(\nX_a1[15] ));
    defparam nX_a1_i15.GSR = "DISABLED";
    FD1S3AX nX_a1_i14 (.D(\nX_a0[14] ), .CK(clock), .Q(\nX_a1[14] ));
    defparam nX_a1_i14.GSR = "DISABLED";
    FD1S3AX nX_a1_i13 (.D(\nX_a0[13] ), .CK(clock), .Q(\nX_a1[13] ));
    defparam nX_a1_i13.GSR = "DISABLED";
    FD1S3AX nX_a1_i12 (.D(\nX_a0[12] ), .CK(clock), .Q(\nX_a1[12] ));
    defparam nX_a1_i12.GSR = "DISABLED";
    FD1S3AX nX_a1_i11 (.D(\nX_a0[11] ), .CK(clock), .Q(\nX_a1[11] ));
    defparam nX_a1_i11.GSR = "DISABLED";
    FD1S3AX nX_a1_i10 (.D(\nX_a0[10] ), .CK(clock), .Q(\nX_a1[10] ));
    defparam nX_a1_i10.GSR = "DISABLED";
    FD1S3AX nX_a1_i9 (.D(\nX_a0[9] ), .CK(clock), .Q(\nX_a1[9] ));
    defparam nX_a1_i9.GSR = "DISABLED";
    FD1S3IX nX_a1_i8 (.D(\buf_x[471] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[8] ));
    defparam nX_a1_i8.GSR = "DISABLED";
    FD1S3IX nX_a1_i7 (.D(\buf_x[470] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[7] ));
    defparam nX_a1_i7.GSR = "DISABLED";
    FD1S3IX nX_a1_i6 (.D(\buf_x[469] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[6] ));
    defparam nX_a1_i6.GSR = "DISABLED";
    FD1S3IX nX_a1_i5 (.D(\buf_x[468] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[5] ));
    defparam nX_a1_i5.GSR = "DISABLED";
    FD1S3IX nX_a1_i4 (.D(\buf_x[467] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[4] ));
    defparam nX_a1_i4.GSR = "DISABLED";
    FD1S3IX nX_a1_i3 (.D(\buf_x[466] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[3] ));
    defparam nX_a1_i3.GSR = "DISABLED";
    FD1S3IX nX_a1_i2 (.D(\buf_x[465] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[2] ));
    defparam nX_a1_i2.GSR = "DISABLED";
    FD1S3IX nX_a1_i1 (.D(\buf_x[464] ), .CK(clock), .CD(\eX_x[11] ), .Q(\nX_a1[1] ));
    defparam nX_a1_i1.GSR = "DISABLED";
    CCU2D add_2948_14 (.A0(buf_x[432]), .B0(buf_x[446]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61737), .S0(\nK0_b0[21] ));
    defparam add_2948_14.INIT0 = 16'h5666;
    defparam add_2948_14.INIT1 = 16'h0000;
    defparam add_2948_14.INJECT1_0 = "NO";
    defparam add_2948_14.INJECT1_1 = "NO";
    CCU2D add_2948_12 (.A0(buf_x[431]), .B0(buf_x[444]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[432]), .B1(buf_x[446]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61736), .COUT(n61737), .S0(\nK0_b0[19] ), 
          .S1(\nK0_b0[20] ));
    defparam add_2948_12.INIT0 = 16'h5666;
    defparam add_2948_12.INIT1 = 16'h5666;
    defparam add_2948_12.INJECT1_0 = "NO";
    defparam add_2948_12.INJECT1_1 = "NO";
    CCU2D add_2948_10 (.A0(buf_x[429]), .B0(buf_x[442]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[430]), .B1(buf_x[443]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61735), .COUT(n61736), .S0(\nK0_b0[17] ), 
          .S1(\nK0_b0[18] ));
    defparam add_2948_10.INIT0 = 16'h5666;
    defparam add_2948_10.INIT1 = 16'h5666;
    defparam add_2948_10.INJECT1_0 = "NO";
    defparam add_2948_10.INJECT1_1 = "NO";
    CCU2D add_2948_8 (.A0(buf_x[427]), .B0(buf_x[440]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[428]), .B1(buf_x[441]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61734), .COUT(n61735), .S0(\nK0_b0[15] ), 
          .S1(\nK0_b0[16] ));
    defparam add_2948_8.INIT0 = 16'h5666;
    defparam add_2948_8.INIT1 = 16'h5666;
    defparam add_2948_8.INJECT1_0 = "NO";
    defparam add_2948_8.INJECT1_1 = "NO";
    CCU2D add_2948_6 (.A0(buf_x[425]), .B0(buf_x[438]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[426]), .B1(buf_x[439]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61733), .COUT(n61734), .S0(\nK0_b0[13] ), 
          .S1(\nK0_b0[14] ));
    defparam add_2948_6.INIT0 = 16'h5666;
    defparam add_2948_6.INIT1 = 16'h5666;
    defparam add_2948_6.INJECT1_0 = "NO";
    defparam add_2948_6.INJECT1_1 = "NO";
    CCU2D add_2948_4 (.A0(buf_x[423]), .B0(\buf_x[436] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[424]), .B1(\buf_x[437] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61732), .COUT(n61733), .S1(\nK0_b0[12] ));
    defparam add_2948_4.INIT0 = 16'h5666;
    defparam add_2948_4.INIT1 = 16'h5666;
    defparam add_2948_4.INJECT1_0 = "NO";
    defparam add_2948_4.INJECT1_1 = "NO";
    CCU2D add_2948_2 (.A0(buf_x[421]), .B0(\buf_x[434] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[422]), .B1(\buf_x[435] ), .C1(GND_net), 
          .D1(GND_net), .COUT(n61732));
    defparam add_2948_2.INIT0 = 16'h7000;
    defparam add_2948_2.INIT1 = 16'h5666;
    defparam add_2948_2.INJECT1_0 = "NO";
    defparam add_2948_2.INJECT1_1 = "NO";
    CCU2D add_19_16 (.A0(buf_x[268]), .B0(buf_x[357]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61731), 
          .S0(buf_x[377]));
    defparam add_19_16.INIT0 = 16'h5666;
    defparam add_19_16.INIT1 = 16'h0000;
    defparam add_19_16.INJECT1_0 = "NO";
    defparam add_19_16.INJECT1_1 = "NO";
    CCU2D add_19_14 (.A0(buf_x[268]), .B0(buf_x[356]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[268]), .B1(buf_x[357]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61730), .COUT(n61731), .S0(buf_x[375]), .S1(buf_x[376]));
    defparam add_19_14.INIT0 = 16'h5666;
    defparam add_19_14.INIT1 = 16'h5666;
    defparam add_19_14.INJECT1_0 = "NO";
    defparam add_19_14.INJECT1_1 = "NO";
    CCU2D add_19_12 (.A0(buf_x[268]), .B0(buf_x[354]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[268]), .B1(buf_x[355]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61729), .COUT(n61730), .S0(buf_x[373]), .S1(buf_x[374]));
    defparam add_19_12.INIT0 = 16'h5666;
    defparam add_19_12.INIT1 = 16'h5666;
    defparam add_19_12.INJECT1_0 = "NO";
    defparam add_19_12.INJECT1_1 = "NO";
    CCU2D add_19_10 (.A0(buf_x[388]), .B0(buf_x[352]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[389]), .B1(buf_x[353]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61728), .COUT(n61729), .S0(buf_x[371]), .S1(buf_x[372]));
    defparam add_19_10.INIT0 = 16'h5666;
    defparam add_19_10.INIT1 = 16'h5666;
    defparam add_19_10.INJECT1_0 = "NO";
    defparam add_19_10.INJECT1_1 = "NO";
    CCU2D add_19_8 (.A0(buf_x[386]), .B0(buf_x[350]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[387]), .B1(buf_x[351]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61727), .COUT(n61728), .S0(buf_x[369]), .S1(buf_x[370]));
    defparam add_19_8.INIT0 = 16'h5666;
    defparam add_19_8.INIT1 = 16'h5666;
    defparam add_19_8.INJECT1_0 = "NO";
    defparam add_19_8.INJECT1_1 = "NO";
    CCU2D add_19_6 (.A0(buf_x[384]), .B0(buf_x[273]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[385]), .B1(buf_x[349]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61726), .COUT(n61727), .S0(buf_x[367]), .S1(buf_x[368]));
    defparam add_19_6.INIT0 = 16'h5666;
    defparam add_19_6.INIT1 = 16'h5666;
    defparam add_19_6.INJECT1_0 = "NO";
    defparam add_19_6.INJECT1_1 = "NO";
    CCU2D add_19_4 (.A0(buf_x[382]), .B0(buf_x[271]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[383]), .B1(buf_x[272]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61725), .COUT(n61726), .S0(buf_x[365]), .S1(buf_x[366]));
    defparam add_19_4.INIT0 = 16'h5666;
    defparam add_19_4.INIT1 = 16'h5666;
    defparam add_19_4.INJECT1_0 = "NO";
    defparam add_19_4.INJECT1_1 = "NO";
    CCU2D add_19_2 (.A0(buf_x[380]), .B0(buf_x[379]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[380]), .B1(buf_x[379]), .C1(buf_x[381]), .D1(GND_net), 
          .COUT(n61725), .S1(buf_x[364]));
    defparam add_19_2.INIT0 = 16'h7000;
    defparam add_19_2.INIT1 = 16'h9696;
    defparam add_19_2.INJECT1_0 = "NO";
    defparam add_19_2.INJECT1_1 = "NO";
    CCU2D add_2947_16 (.A0(buf_r[357]), .B0(buf_r[376]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[357]), .B1(buf_r[377]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61722), .S0(buf_x[431]), .S1(buf_x[432]));
    defparam add_2947_16.INIT0 = 16'h5666;
    defparam add_2947_16.INIT1 = 16'h5666;
    defparam add_2947_16.INJECT1_0 = "NO";
    defparam add_2947_16.INJECT1_1 = "NO";
    CCU2D add_2947_14 (.A0(buf_r[357]), .B0(buf_r[374]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[357]), .B1(buf_r[375]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61721), .COUT(n61722), .S0(buf_x[429]), 
          .S1(buf_x[430]));
    defparam add_2947_14.INIT0 = 16'h5666;
    defparam add_2947_14.INIT1 = 16'h5666;
    defparam add_2947_14.INJECT1_0 = "NO";
    defparam add_2947_14.INJECT1_1 = "NO";
    CCU2D add_2947_12 (.A0(buf_r[357]), .B0(buf_r[372]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[357]), .B1(buf_r[373]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61720), .COUT(n61721), .S0(buf_x[427]), 
          .S1(buf_x[428]));
    defparam add_2947_12.INIT0 = 16'h5666;
    defparam add_2947_12.INIT1 = 16'h5666;
    defparam add_2947_12.INJECT1_0 = "NO";
    defparam add_2947_12.INJECT1_1 = "NO";
    CCU2D add_2947_10 (.A0(buf_r[357]), .B0(buf_r[370]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[357]), .B1(buf_r[371]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61719), .COUT(n61720), .S0(buf_x[425]), 
          .S1(buf_x[426]));
    defparam add_2947_10.INIT0 = 16'h5666;
    defparam add_2947_10.INIT1 = 16'h5666;
    defparam add_2947_10.INJECT1_0 = "NO";
    defparam add_2947_10.INJECT1_1 = "NO";
    CCU2D add_2947_8 (.A0(buf_r[355]), .B0(buf_r[368]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[356]), .B1(buf_r[369]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61718), .COUT(n61719), .S0(buf_x[423]), 
          .S1(buf_x[424]));
    defparam add_2947_8.INIT0 = 16'h5666;
    defparam add_2947_8.INIT1 = 16'h5666;
    defparam add_2947_8.INJECT1_0 = "NO";
    defparam add_2947_8.INJECT1_1 = "NO";
    CCU2D add_2947_6 (.A0(buf_r[353]), .B0(buf_r[366]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[354]), .B1(buf_r[367]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61717), .COUT(n61718), .S0(buf_x[421]), 
          .S1(buf_x[422]));
    defparam add_2947_6.INIT0 = 16'h5666;
    defparam add_2947_6.INIT1 = 16'h5666;
    defparam add_2947_6.INJECT1_0 = "NO";
    defparam add_2947_6.INJECT1_1 = "NO";
    CCU2D add_2947_4 (.A0(buf_r[351]), .B0(buf_r[364]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[352]), .B1(buf_r[365]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61716), .COUT(n61717));
    defparam add_2947_4.INIT0 = 16'h5666;
    defparam add_2947_4.INIT1 = 16'h5666;
    defparam add_2947_4.INJECT1_0 = "NO";
    defparam add_2947_4.INJECT1_1 = "NO";
    CCU2D add_2947_2 (.A0(buf_r[349]), .B0(\buf_x[434] ), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[350]), .B1(buf_r[363]), .C1(GND_net), 
          .D1(GND_net), .COUT(n61716));
    defparam add_2947_2.INIT0 = 16'h7000;
    defparam add_2947_2.INIT1 = 16'h5666;
    defparam add_2947_2.INJECT1_0 = "NO";
    defparam add_2947_2.INJECT1_1 = "NO";
    CCU2D add_16_14 (.A0(buf_x[268]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61715), 
          .S0(buf_x[357]));
    defparam add_16_14.INIT0 = 16'h5000;
    defparam add_16_14.INIT1 = 16'h0000;
    defparam add_16_14.INJECT1_0 = "NO";
    defparam add_16_14.INJECT1_1 = "NO";
    CCU2D add_16_12 (.A0(buf_x[268]), .B0(buf_x[389]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[268]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61714), .COUT(n61715), .S0(buf_x[355]), .S1(buf_x[356]));
    defparam add_16_12.INIT0 = 16'h5666;
    defparam add_16_12.INIT1 = 16'h5000;
    defparam add_16_12.INJECT1_0 = "NO";
    defparam add_16_12.INJECT1_1 = "NO";
    CCU2D add_16_10 (.A0(buf_x[388]), .B0(buf_x[387]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[389]), .B1(buf_x[388]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61713), .COUT(n61714), .S0(buf_x[353]), .S1(buf_x[354]));
    defparam add_16_10.INIT0 = 16'h5666;
    defparam add_16_10.INIT1 = 16'h5666;
    defparam add_16_10.INJECT1_0 = "NO";
    defparam add_16_10.INJECT1_1 = "NO";
    CCU2D add_16_8 (.A0(buf_x[386]), .B0(buf_x[385]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[387]), .B1(buf_x[386]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61712), .COUT(n61713), .S0(buf_x[351]), .S1(buf_x[352]));
    defparam add_16_8.INIT0 = 16'h5666;
    defparam add_16_8.INIT1 = 16'h5666;
    defparam add_16_8.INJECT1_0 = "NO";
    defparam add_16_8.INJECT1_1 = "NO";
    CCU2D add_16_6 (.A0(buf_x[384]), .B0(buf_x[383]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[385]), .B1(buf_x[384]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61711), .COUT(n61712), .S0(buf_x[349]), .S1(buf_x[350]));
    defparam add_16_6.INIT0 = 16'h5666;
    defparam add_16_6.INIT1 = 16'h5666;
    defparam add_16_6.INJECT1_0 = "NO";
    defparam add_16_6.INJECT1_1 = "NO";
    CCU2D add_16_4 (.A0(buf_x[382]), .B0(buf_x[381]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[383]), .B1(buf_x[382]), .C1(GND_net), .D1(GND_net), 
          .CIN(n61710), .COUT(n61711), .S0(buf_x[272]), .S1(buf_x[273]));
    defparam add_16_4.INIT0 = 16'h5666;
    defparam add_16_4.INIT1 = 16'h5666;
    defparam add_16_4.INJECT1_0 = "NO";
    defparam add_16_4.INJECT1_1 = "NO";
    CCU2D add_16_2 (.A0(buf_x[380]), .B0(buf_x[379]), .C0(GND_net), .D0(GND_net), 
          .A1(buf_x[381]), .B1(buf_x[380]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61710), .S1(buf_x[271]));
    defparam add_16_2.INIT0 = 16'h7000;
    defparam add_16_2.INIT1 = 16'h5666;
    defparam add_16_2.INJECT1_0 = "NO";
    defparam add_16_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \fp_exp_exp_y2_clk(23) 
//

module \fp_exp_exp_y2_clk(23)  (\buf[50] , \buf[51] , \buf[52] , \buf[53] , 
            \buf[54] , \buf[55] , \r_0[6] , \r_0[7] , \r_0[8] , n15447, 
            n15462, GND_net, nEY2_d1, n15449, n15448, n15451, n15450, 
            n15453, n15469, n15452, n15455, n15471, n15454, n15470, 
            n15457, n15473, n15456, n15472, n15459, n15475, n15458, 
            n15474, \nY_c1[8] , \nY_c1[13] , \r_1[7] , clock, \r_1[6] , 
            \r_1[5] , \r_1[4] , \r_1[3] , \r_1[2] , \r_1[1] , \r_1[0] , 
            \nY_c1[20] , \nY_c1[21] , \nY_c1[22] , \nY_c1[23] , \nY_c1[24] , 
            \nY_c1[25] , \nY_c1[26] , \nY1_c1[7] , \nEY1_c1[9] , \nEY1_c1[10] , 
            \nEY1_c1[11] , \nEY1_c1[12] , \nEY1_c1[13] , \nEY1_c1[14] , 
            \nEY1_c1[15] , \nEY1_c1[16] , \nEY1_c1[17] , \nEY1_c1[0] , 
            \nEY1_c1[1] , \nEY1_c1[2] , \nEY1_c1[3] , \nEY1_c1[4] , 
            \nEY1_c1[5] , \nEY1_c1[6] , \nEY1_c1[7] , \nEY1_c1[8] , 
            VCC_net, \nY_c1[10] , \nY_c1[12] , \nEY1_c1[19] , \nEY1_c1[20] , 
            \nEY1_c1[21] , \nEY1_c1[22] , \nEY1_c1[23] , \nEY1_c1[24] , 
            \nEY1_c1[18] , \nY_c1[19] , \nY_c1[18] , \nY_c1[17] , \nY_c1[16] , 
            \nY_c1[15] , \nY_c1[14] , \nY_c1[11] , \nY_c1[9] , \buf_x[89] , 
            \buf_x[87] , \buf_x[88] , \buf_x[85] , \buf_x[86] , \buf_x[83] , 
            \buf_x[84] , \buf_r[89] , \buf_r[87] , \buf_r[88] , \buf_r[85] , 
            \buf_r[86] , \buf_r[83] , \buf_r[84] );
    input \buf[50] ;
    input \buf[51] ;
    input \buf[52] ;
    input \buf[53] ;
    input \buf[54] ;
    input \buf[55] ;
    output \r_0[6] ;
    output \r_0[7] ;
    output \r_0[8] ;
    input n15447;
    input n15462;
    input GND_net;
    output [12:0]nEY2_d1;
    input n15449;
    input n15448;
    input n15451;
    input n15450;
    input n15453;
    input n15469;
    input n15452;
    input n15455;
    input n15471;
    input n15454;
    input n15470;
    input n15457;
    input n15473;
    input n15456;
    input n15472;
    input n15459;
    input n15475;
    input n15458;
    input n15474;
    input \nY_c1[8] ;
    input \nY_c1[13] ;
    output \r_1[7] ;
    input clock;
    output \r_1[6] ;
    output \r_1[5] ;
    output \r_1[4] ;
    output \r_1[3] ;
    output \r_1[2] ;
    output \r_1[1] ;
    output \r_1[0] ;
    input \nY_c1[20] ;
    input \nY_c1[21] ;
    input \nY_c1[22] ;
    input \nY_c1[23] ;
    input \nY_c1[24] ;
    input \nY_c1[25] ;
    input \nY_c1[26] ;
    input \nY1_c1[7] ;
    output \nEY1_c1[9] ;
    output \nEY1_c1[10] ;
    output \nEY1_c1[11] ;
    output \nEY1_c1[12] ;
    output \nEY1_c1[13] ;
    output \nEY1_c1[14] ;
    output \nEY1_c1[15] ;
    output \nEY1_c1[16] ;
    output \nEY1_c1[17] ;
    output \nEY1_c1[0] ;
    output \nEY1_c1[1] ;
    output \nEY1_c1[2] ;
    output \nEY1_c1[3] ;
    output \nEY1_c1[4] ;
    output \nEY1_c1[5] ;
    output \nEY1_c1[6] ;
    output \nEY1_c1[7] ;
    output \nEY1_c1[8] ;
    input VCC_net;
    input \nY_c1[10] ;
    input \nY_c1[12] ;
    output \nEY1_c1[19] ;
    output \nEY1_c1[20] ;
    output \nEY1_c1[21] ;
    output \nEY1_c1[22] ;
    output \nEY1_c1[23] ;
    output \nEY1_c1[24] ;
    output \nEY1_c1[18] ;
    input \nY_c1[19] ;
    input \nY_c1[18] ;
    input \nY_c1[17] ;
    input \nY_c1[16] ;
    input \nY_c1[15] ;
    input \nY_c1[14] ;
    input \nY_c1[11] ;
    input \nY_c1[9] ;
    output \buf_x[89] ;
    output \buf_x[87] ;
    output \buf_x[88] ;
    output \buf_x[85] ;
    output \buf_x[86] ;
    output \buf_x[83] ;
    output \buf_x[84] ;
    input \buf_r[89] ;
    input \buf_r[87] ;
    input \buf_r[88] ;
    input \buf_r[85] ;
    input \buf_r[86] ;
    input \buf_r[83] ;
    input \buf_r[84] ;
    
    
    fp_exp_exp_y2_23_clk \exp_y2_23.exp_y2  (.\buf[50] (\buf[50] ), .\buf[51] (\buf[51] ), 
            .\buf[52] (\buf[52] ), .\buf[53] (\buf[53] ), .\buf[54] (\buf[54] ), 
            .\buf[55] (\buf[55] ), .\r_0[6] (\r_0[6] ), .\r_0[7] (\r_0[7] ), 
            .\r_0[8] (\r_0[8] ), .n15447(n15447), .n15462(n15462), .GND_net(GND_net), 
            .nEY2_d1({nEY2_d1}), .n15449(n15449), .n15448(n15448), .n15451(n15451), 
            .n15450(n15450), .n15453(n15453), .n15469(n15469), .n15452(n15452), 
            .n15455(n15455), .n15471(n15471), .n15454(n15454), .n15470(n15470), 
            .n15457(n15457), .n15473(n15473), .n15456(n15456), .n15472(n15472), 
            .n15459(n15459), .n15475(n15475), .n15458(n15458), .n15474(n15474), 
            .\nY_c1[8] (\nY_c1[8] ), .\nY_c1[13] (\nY_c1[13] ), .\r_1[7] (\r_1[7] ), 
            .clock(clock), .\r_1[6] (\r_1[6] ), .\r_1[5] (\r_1[5] ), .\r_1[4] (\r_1[4] ), 
            .\r_1[3] (\r_1[3] ), .\r_1[2] (\r_1[2] ), .\r_1[1] (\r_1[1] ), 
            .\r_1[0] (\r_1[0] ), .\nY_c1[20] (\nY_c1[20] ), .\nY_c1[21] (\nY_c1[21] ), 
            .\nY_c1[22] (\nY_c1[22] ), .\nY_c1[23] (\nY_c1[23] ), .\nY_c1[24] (\nY_c1[24] ), 
            .\nY_c1[25] (\nY_c1[25] ), .\nY_c1[26] (\nY_c1[26] ), .\nY1_c1[7] (\nY1_c1[7] ), 
            .\nEY1_c1[9] (\nEY1_c1[9] ), .\nEY1_c1[10] (\nEY1_c1[10] ), 
            .\nEY1_c1[11] (\nEY1_c1[11] ), .\nEY1_c1[12] (\nEY1_c1[12] ), 
            .\nEY1_c1[13] (\nEY1_c1[13] ), .\nEY1_c1[14] (\nEY1_c1[14] ), 
            .\nEY1_c1[15] (\nEY1_c1[15] ), .\nEY1_c1[16] (\nEY1_c1[16] ), 
            .\nEY1_c1[17] (\nEY1_c1[17] ), .\nEY1_c1[0] (\nEY1_c1[0] ), 
            .\nEY1_c1[1] (\nEY1_c1[1] ), .\nEY1_c1[2] (\nEY1_c1[2] ), .\nEY1_c1[3] (\nEY1_c1[3] ), 
            .\nEY1_c1[4] (\nEY1_c1[4] ), .\nEY1_c1[5] (\nEY1_c1[5] ), .\nEY1_c1[6] (\nEY1_c1[6] ), 
            .\nEY1_c1[7] (\nEY1_c1[7] ), .\nEY1_c1[8] (\nEY1_c1[8] ), .VCC_net(VCC_net), 
            .\nY_c1[10] (\nY_c1[10] ), .\nY_c1[12] (\nY_c1[12] ), .\nEY1_c1[19] (\nEY1_c1[19] ), 
            .\nEY1_c1[20] (\nEY1_c1[20] ), .\nEY1_c1[21] (\nEY1_c1[21] ), 
            .\nEY1_c1[22] (\nEY1_c1[22] ), .\nEY1_c1[23] (\nEY1_c1[23] ), 
            .\nEY1_c1[24] (\nEY1_c1[24] ), .\nEY1_c1[18] (\nEY1_c1[18] ), 
            .\nY_c1[19] (\nY_c1[19] ), .\nY_c1[18] (\nY_c1[18] ), .\nY_c1[17] (\nY_c1[17] ), 
            .\nY_c1[16] (\nY_c1[16] ), .\nY_c1[15] (\nY_c1[15] ), .\nY_c1[14] (\nY_c1[14] ), 
            .\nY_c1[11] (\nY_c1[11] ), .\nY_c1[9] (\nY_c1[9] ), .\buf_x[89] (\buf_x[89] ), 
            .\buf_x[87] (\buf_x[87] ), .\buf_x[88] (\buf_x[88] ), .\buf_x[85] (\buf_x[85] ), 
            .\buf_x[86] (\buf_x[86] ), .\buf_x[83] (\buf_x[83] ), .\buf_x[84] (\buf_x[84] ), 
            .\buf_r[89] (\buf_r[89] ), .\buf_r[87] (\buf_r[87] ), .\buf_r[88] (\buf_r[88] ), 
            .\buf_r[85] (\buf_r[85] ), .\buf_r[86] (\buf_r[86] ), .\buf_r[83] (\buf_r[83] ), 
            .\buf_r[84] (\buf_r[84] ));
    
endmodule
//
// Verilog Description of module fp_exp_exp_y2_23_clk
//

module fp_exp_exp_y2_23_clk (\buf[50] , \buf[51] , \buf[52] , \buf[53] , 
            \buf[54] , \buf[55] , \r_0[6] , \r_0[7] , \r_0[8] , n15447, 
            n15462, GND_net, nEY2_d1, n15449, n15448, n15451, n15450, 
            n15453, n15469, n15452, n15455, n15471, n15454, n15470, 
            n15457, n15473, n15456, n15472, n15459, n15475, n15458, 
            n15474, \nY_c1[8] , \nY_c1[13] , \r_1[7] , clock, \r_1[6] , 
            \r_1[5] , \r_1[4] , \r_1[3] , \r_1[2] , \r_1[1] , \r_1[0] , 
            \nY_c1[20] , \nY_c1[21] , \nY_c1[22] , \nY_c1[23] , \nY_c1[24] , 
            \nY_c1[25] , \nY_c1[26] , \nY1_c1[7] , \nEY1_c1[9] , \nEY1_c1[10] , 
            \nEY1_c1[11] , \nEY1_c1[12] , \nEY1_c1[13] , \nEY1_c1[14] , 
            \nEY1_c1[15] , \nEY1_c1[16] , \nEY1_c1[17] , \nEY1_c1[0] , 
            \nEY1_c1[1] , \nEY1_c1[2] , \nEY1_c1[3] , \nEY1_c1[4] , 
            \nEY1_c1[5] , \nEY1_c1[6] , \nEY1_c1[7] , \nEY1_c1[8] , 
            VCC_net, \nY_c1[10] , \nY_c1[12] , \nEY1_c1[19] , \nEY1_c1[20] , 
            \nEY1_c1[21] , \nEY1_c1[22] , \nEY1_c1[23] , \nEY1_c1[24] , 
            \nEY1_c1[18] , \nY_c1[19] , \nY_c1[18] , \nY_c1[17] , \nY_c1[16] , 
            \nY_c1[15] , \nY_c1[14] , \nY_c1[11] , \nY_c1[9] , \buf_x[89] , 
            \buf_x[87] , \buf_x[88] , \buf_x[85] , \buf_x[86] , \buf_x[83] , 
            \buf_x[84] , \buf_r[89] , \buf_r[87] , \buf_r[88] , \buf_r[85] , 
            \buf_r[86] , \buf_r[83] , \buf_r[84] );
    input \buf[50] ;
    input \buf[51] ;
    input \buf[52] ;
    input \buf[53] ;
    input \buf[54] ;
    input \buf[55] ;
    output \r_0[6] ;
    output \r_0[7] ;
    output \r_0[8] ;
    input n15447;
    input n15462;
    input GND_net;
    output [12:0]nEY2_d1;
    input n15449;
    input n15448;
    input n15451;
    input n15450;
    input n15453;
    input n15469;
    input n15452;
    input n15455;
    input n15471;
    input n15454;
    input n15470;
    input n15457;
    input n15473;
    input n15456;
    input n15472;
    input n15459;
    input n15475;
    input n15458;
    input n15474;
    input \nY_c1[8] ;
    input \nY_c1[13] ;
    output \r_1[7] ;
    input clock;
    output \r_1[6] ;
    output \r_1[5] ;
    output \r_1[4] ;
    output \r_1[3] ;
    output \r_1[2] ;
    output \r_1[1] ;
    output \r_1[0] ;
    input \nY_c1[20] ;
    input \nY_c1[21] ;
    input \nY_c1[22] ;
    input \nY_c1[23] ;
    input \nY_c1[24] ;
    input \nY_c1[25] ;
    input \nY_c1[26] ;
    input \nY1_c1[7] ;
    output \nEY1_c1[9] ;
    output \nEY1_c1[10] ;
    output \nEY1_c1[11] ;
    output \nEY1_c1[12] ;
    output \nEY1_c1[13] ;
    output \nEY1_c1[14] ;
    output \nEY1_c1[15] ;
    output \nEY1_c1[16] ;
    output \nEY1_c1[17] ;
    output \nEY1_c1[0] ;
    output \nEY1_c1[1] ;
    output \nEY1_c1[2] ;
    output \nEY1_c1[3] ;
    output \nEY1_c1[4] ;
    output \nEY1_c1[5] ;
    output \nEY1_c1[6] ;
    output \nEY1_c1[7] ;
    output \nEY1_c1[8] ;
    input VCC_net;
    input \nY_c1[10] ;
    input \nY_c1[12] ;
    output \nEY1_c1[19] ;
    output \nEY1_c1[20] ;
    output \nEY1_c1[21] ;
    output \nEY1_c1[22] ;
    output \nEY1_c1[23] ;
    output \nEY1_c1[24] ;
    output \nEY1_c1[18] ;
    input \nY_c1[19] ;
    input \nY_c1[18] ;
    input \nY_c1[17] ;
    input \nY_c1[16] ;
    input \nY_c1[15] ;
    input \nY_c1[14] ;
    input \nY_c1[11] ;
    input \nY_c1[9] ;
    output \buf_x[89] ;
    output \buf_x[87] ;
    output \buf_x[88] ;
    output \buf_x[85] ;
    output \buf_x[86] ;
    output \buf_x[83] ;
    output \buf_x[84] ;
    input \buf_r[89] ;
    input \buf_r[87] ;
    input \buf_r[88] ;
    input \buf_r[85] ;
    input \buf_r[86] ;
    input \buf_r[83] ;
    input \buf_r[84] ;
    
    
    wire n62195, n62194, n62193, n62192, n62191, n62190;
    
    ROM64X1A Mux_9 (.AD0(\buf[50] ), .AD1(\buf[51] ), .AD2(\buf[52] ), 
            .AD3(\buf[53] ), .AD4(\buf[54] ), .AD5(\buf[55] ), .DO0(\r_0[6] )) /* synthesis initstate=0x07255B3FFCDAA4C0 */ ;
    defparam Mux_9.initval = 64'h07255B3FFCDAA4C0;
    ROM64X1A Mux_8 (.AD0(\buf[50] ), .AD1(\buf[51] ), .AD2(\buf[52] ), 
            .AD3(\buf[53] ), .AD4(\buf[54] ), .AD5(\buf[55] ), .DO0(\r_0[7] )) /* synthesis initstate=0xFF1CC96AA96CC700 */ ;
    defparam Mux_8.initval = 64'hFF1CC96AA96CC700;
    ROM64X1A Mux_7 (.AD0(\buf[50] ), .AD1(\buf[51] ), .AD2(\buf[52] ), 
            .AD3(\buf[53] ), .AD4(\buf[54] ), .AD5(\buf[55] ), .DO0(\r_0[8] )) /* synthesis initstate=0xAA56924CCE70F800 */ ;
    defparam Mux_7.initval = 64'hAA56924CCE70F800;
    CCU2D add_4_14 (.A0(n15447), .B0(n15462), .C0(GND_net), .D0(GND_net), 
          .A1(n15462), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62195), 
          .S0(nEY2_d1[11]), .S1(nEY2_d1[12]));
    defparam add_4_14.INIT0 = 16'h5666;
    defparam add_4_14.INIT1 = 16'hfaaa;
    defparam add_4_14.INJECT1_0 = "NO";
    defparam add_4_14.INJECT1_1 = "NO";
    CCU2D add_4_12 (.A0(n15449), .B0(n15462), .C0(GND_net), .D0(GND_net), 
          .A1(n15448), .B1(n15462), .C1(GND_net), .D1(GND_net), .CIN(n62194), 
          .COUT(n62195), .S0(nEY2_d1[9]), .S1(nEY2_d1[10]));
    defparam add_4_12.INIT0 = 16'h5666;
    defparam add_4_12.INIT1 = 16'h5666;
    defparam add_4_12.INJECT1_0 = "NO";
    defparam add_4_12.INJECT1_1 = "NO";
    CCU2D add_4_10 (.A0(n15451), .B0(n15462), .C0(GND_net), .D0(GND_net), 
          .A1(n15450), .B1(n15462), .C1(GND_net), .D1(GND_net), .CIN(n62193), 
          .COUT(n62194), .S0(nEY2_d1[7]), .S1(nEY2_d1[8]));
    defparam add_4_10.INIT0 = 16'h5666;
    defparam add_4_10.INIT1 = 16'h5666;
    defparam add_4_10.INJECT1_0 = "NO";
    defparam add_4_10.INJECT1_1 = "NO";
    CCU2D add_4_8 (.A0(n15453), .B0(n15469), .C0(GND_net), .D0(GND_net), 
          .A1(n15452), .B1(n15462), .C1(GND_net), .D1(GND_net), .CIN(n62192), 
          .COUT(n62193), .S0(nEY2_d1[5]), .S1(nEY2_d1[6]));
    defparam add_4_8.INIT0 = 16'h5666;
    defparam add_4_8.INIT1 = 16'h5666;
    defparam add_4_8.INJECT1_0 = "NO";
    defparam add_4_8.INJECT1_1 = "NO";
    CCU2D add_4_6 (.A0(n15455), .B0(n15471), .C0(GND_net), .D0(GND_net), 
          .A1(n15454), .B1(n15470), .C1(GND_net), .D1(GND_net), .CIN(n62191), 
          .COUT(n62192), .S0(nEY2_d1[3]), .S1(nEY2_d1[4]));
    defparam add_4_6.INIT0 = 16'h5666;
    defparam add_4_6.INIT1 = 16'h5666;
    defparam add_4_6.INJECT1_0 = "NO";
    defparam add_4_6.INJECT1_1 = "NO";
    CCU2D add_4_4 (.A0(n15457), .B0(n15473), .C0(GND_net), .D0(GND_net), 
          .A1(n15456), .B1(n15472), .C1(GND_net), .D1(GND_net), .CIN(n62190), 
          .COUT(n62191), .S0(nEY2_d1[1]), .S1(nEY2_d1[2]));
    defparam add_4_4.INIT0 = 16'h5666;
    defparam add_4_4.INIT1 = 16'h5666;
    defparam add_4_4.INJECT1_0 = "NO";
    defparam add_4_4.INJECT1_1 = "NO";
    CCU2D add_4_2 (.A0(n15459), .B0(n15475), .C0(GND_net), .D0(GND_net), 
          .A1(n15458), .B1(n15474), .C1(GND_net), .D1(GND_net), .COUT(n62190), 
          .S1(nEY2_d1[0]));
    defparam add_4_2.INIT0 = 16'h7000;
    defparam add_4_2.INIT1 = 16'h5666;
    defparam add_4_2.INJECT1_0 = "NO";
    defparam add_4_2.INJECT1_1 = "NO";
    fp_exp_exp_y2_23_t1_clk t_1 (.\nY_c1[8] (\nY_c1[8] ), .\nY_c1[13] (\nY_c1[13] ), 
            .\r_1[7] (\r_1[7] ), .clock(clock), .\r_1[6] (\r_1[6] ), .\r_1[5] (\r_1[5] ), 
            .\r_1[4] (\r_1[4] ), .\r_1[3] (\r_1[3] ), .\r_1[2] (\r_1[2] ), 
            .\r_1[1] (\r_1[1] ), .\r_1[0] (\r_1[0] ), .\nY_c1[20] (\nY_c1[20] ), 
            .\nY_c1[21] (\nY_c1[21] ), .\nY_c1[22] (\nY_c1[22] ), .\nY_c1[23] (\nY_c1[23] ), 
            .\nY_c1[24] (\nY_c1[24] ), .\nY_c1[25] (\nY_c1[25] ), .\nY_c1[26] (\nY_c1[26] ), 
            .\nY1_c1[7] (\nY1_c1[7] ), .\nEY1_c1[9] (\nEY1_c1[9] ), .\nEY1_c1[10] (\nEY1_c1[10] ), 
            .\nEY1_c1[11] (\nEY1_c1[11] ), .\nEY1_c1[12] (\nEY1_c1[12] ), 
            .\nEY1_c1[13] (\nEY1_c1[13] ), .\nEY1_c1[14] (\nEY1_c1[14] ), 
            .\nEY1_c1[15] (\nEY1_c1[15] ), .\nEY1_c1[16] (\nEY1_c1[16] ), 
            .\nEY1_c1[17] (\nEY1_c1[17] ), .\nEY1_c1[0] (\nEY1_c1[0] ), 
            .\nEY1_c1[1] (\nEY1_c1[1] ), .\nEY1_c1[2] (\nEY1_c1[2] ), .\nEY1_c1[3] (\nEY1_c1[3] ), 
            .\nEY1_c1[4] (\nEY1_c1[4] ), .\nEY1_c1[5] (\nEY1_c1[5] ), .\nEY1_c1[6] (\nEY1_c1[6] ), 
            .\nEY1_c1[7] (\nEY1_c1[7] ), .\nEY1_c1[8] (\nEY1_c1[8] ), .GND_net(GND_net), 
            .VCC_net(VCC_net), .\nY_c1[10] (\nY_c1[10] ), .\nY_c1[12] (\nY_c1[12] ), 
            .\nEY1_c1[19] (\nEY1_c1[19] ), .\nEY1_c1[20] (\nEY1_c1[20] ), 
            .\nEY1_c1[21] (\nEY1_c1[21] ), .\nEY1_c1[22] (\nEY1_c1[22] ), 
            .\nEY1_c1[23] (\nEY1_c1[23] ), .\nEY1_c1[24] (\nEY1_c1[24] ), 
            .\nEY1_c1[18] (\nEY1_c1[18] ), .\nY_c1[19] (\nY_c1[19] ), .\nY_c1[18] (\nY_c1[18] ), 
            .\nY_c1[17] (\nY_c1[17] ), .\nY_c1[16] (\nY_c1[16] ), .\nY_c1[15] (\nY_c1[15] ), 
            .\nY_c1[14] (\nY_c1[14] ), .\nY_c1[11] (\nY_c1[11] ), .\nY_c1[9] (\nY_c1[9] ), 
            .\buf_x[89] (\buf_x[89] ), .\buf_x[87] (\buf_x[87] ), .\buf_x[88] (\buf_x[88] ), 
            .\buf_x[85] (\buf_x[85] ), .\buf_x[86] (\buf_x[86] ), .\buf_x[83] (\buf_x[83] ), 
            .\buf_x[84] (\buf_x[84] ), .\buf_r[89] (\buf_r[89] ), .\buf_r[87] (\buf_r[87] ), 
            .\buf_r[88] (\buf_r[88] ), .\buf_r[85] (\buf_r[85] ), .\buf_r[86] (\buf_r[86] ), 
            .\buf_r[83] (\buf_r[83] ), .\buf_r[84] (\buf_r[84] ));
    
endmodule
//
// Verilog Description of module fp_exp_exp_y2_23_t1_clk
//

module fp_exp_exp_y2_23_t1_clk (\nY_c1[8] , \nY_c1[13] , \r_1[7] , clock, 
            \r_1[6] , \r_1[5] , \r_1[4] , \r_1[3] , \r_1[2] , \r_1[1] , 
            \r_1[0] , \nY_c1[20] , \nY_c1[21] , \nY_c1[22] , \nY_c1[23] , 
            \nY_c1[24] , \nY_c1[25] , \nY_c1[26] , \nY1_c1[7] , \nEY1_c1[9] , 
            \nEY1_c1[10] , \nEY1_c1[11] , \nEY1_c1[12] , \nEY1_c1[13] , 
            \nEY1_c1[14] , \nEY1_c1[15] , \nEY1_c1[16] , \nEY1_c1[17] , 
            \nEY1_c1[0] , \nEY1_c1[1] , \nEY1_c1[2] , \nEY1_c1[3] , 
            \nEY1_c1[4] , \nEY1_c1[5] , \nEY1_c1[6] , \nEY1_c1[7] , 
            \nEY1_c1[8] , GND_net, VCC_net, \nY_c1[10] , \nY_c1[12] , 
            \nEY1_c1[19] , \nEY1_c1[20] , \nEY1_c1[21] , \nEY1_c1[22] , 
            \nEY1_c1[23] , \nEY1_c1[24] , \nEY1_c1[18] , \nY_c1[19] , 
            \nY_c1[18] , \nY_c1[17] , \nY_c1[16] , \nY_c1[15] , \nY_c1[14] , 
            \nY_c1[11] , \nY_c1[9] , \buf_x[89] , \buf_x[87] , \buf_x[88] , 
            \buf_x[85] , \buf_x[86] , \buf_x[83] , \buf_x[84] , \buf_r[89] , 
            \buf_r[87] , \buf_r[88] , \buf_r[85] , \buf_r[86] , \buf_r[83] , 
            \buf_r[84] );
    input \nY_c1[8] ;
    input \nY_c1[13] ;
    output \r_1[7] ;
    input clock;
    output \r_1[6] ;
    output \r_1[5] ;
    output \r_1[4] ;
    output \r_1[3] ;
    output \r_1[2] ;
    output \r_1[1] ;
    output \r_1[0] ;
    input \nY_c1[20] ;
    input \nY_c1[21] ;
    input \nY_c1[22] ;
    input \nY_c1[23] ;
    input \nY_c1[24] ;
    input \nY_c1[25] ;
    input \nY_c1[26] ;
    input \nY1_c1[7] ;
    output \nEY1_c1[9] ;
    output \nEY1_c1[10] ;
    output \nEY1_c1[11] ;
    output \nEY1_c1[12] ;
    output \nEY1_c1[13] ;
    output \nEY1_c1[14] ;
    output \nEY1_c1[15] ;
    output \nEY1_c1[16] ;
    output \nEY1_c1[17] ;
    output \nEY1_c1[0] ;
    output \nEY1_c1[1] ;
    output \nEY1_c1[2] ;
    output \nEY1_c1[3] ;
    output \nEY1_c1[4] ;
    output \nEY1_c1[5] ;
    output \nEY1_c1[6] ;
    output \nEY1_c1[7] ;
    output \nEY1_c1[8] ;
    input GND_net;
    input VCC_net;
    input \nY_c1[10] ;
    input \nY_c1[12] ;
    output \nEY1_c1[19] ;
    output \nEY1_c1[20] ;
    output \nEY1_c1[21] ;
    output \nEY1_c1[22] ;
    output \nEY1_c1[23] ;
    output \nEY1_c1[24] ;
    output \nEY1_c1[18] ;
    input \nY_c1[19] ;
    input \nY_c1[18] ;
    input \nY_c1[17] ;
    input \nY_c1[16] ;
    input \nY_c1[15] ;
    input \nY_c1[14] ;
    input \nY_c1[11] ;
    input \nY_c1[9] ;
    output \buf_x[89] ;
    output \buf_x[87] ;
    output \buf_x[88] ;
    output \buf_x[85] ;
    output \buf_x[86] ;
    output \buf_x[83] ;
    output \buf_x[84] ;
    input \buf_r[89] ;
    input \buf_r[87] ;
    input \buf_r[88] ;
    input \buf_r[85] ;
    input \buf_r[86] ;
    input \buf_r[83] ;
    input \buf_r[84] ;
    
    wire [5:0]s_1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(7594[10:13])
    wire sign_x0;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(7598[10:17])
    wire [14:0]r0_1;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(7596[10:14])
    
    wire n70818;
    
    LUT4 i10013_1_lut_2_lut (.A(\nY_c1[8] ), .B(\nY_c1[13] ), .Z(s_1[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i10013_1_lut_2_lut.init = 16'h9999;
    LUT4 i1_2_lut_rep_848 (.A(\nY_c1[8] ), .B(\nY_c1[13] ), .Z(n70818)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_848.init = 16'h6666;
    FD1S3AX sign_xr_11 (.D(sign_x0), .CK(clock), .Q(\r_1[7] ));
    defparam sign_xr_11.GSR = "DISABLED";
    LUT4 i4_1_lut (.A(\nY_c1[13] ), .Z(sign_x0)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4_1_lut.init = 16'h5555;
    LUT4 xor_9_i7_2_lut (.A(r0_1[13]), .B(\r_1[7] ), .Z(\r_1[6] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i7_2_lut.init = 16'h6666;
    LUT4 xor_9_i6_2_lut (.A(r0_1[12]), .B(\r_1[7] ), .Z(\r_1[5] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i6_2_lut.init = 16'h6666;
    LUT4 xor_9_i5_2_lut (.A(r0_1[11]), .B(\r_1[7] ), .Z(\r_1[4] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i5_2_lut.init = 16'h6666;
    LUT4 xor_9_i4_2_lut (.A(r0_1[10]), .B(\r_1[7] ), .Z(\r_1[3] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i4_2_lut.init = 16'h6666;
    LUT4 xor_9_i3_2_lut (.A(r0_1[9]), .B(\r_1[7] ), .Z(\r_1[2] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i3_2_lut.init = 16'h6666;
    LUT4 xor_9_i2_2_lut (.A(r0_1[8]), .B(\r_1[7] ), .Z(\r_1[1] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i2_2_lut.init = 16'h6666;
    LUT4 xor_9_i1_2_lut (.A(r0_1[7]), .B(\r_1[7] ), .Z(\r_1[0] )) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam xor_9_i1_2_lut.init = 16'h6666;
    \mult_clk(8,6,false,false,1,3)  mult_r0_1 (.\nY_c1[20] (\nY_c1[20] ), 
            .\nY_c1[21] (\nY_c1[21] ), .\nY_c1[22] (\nY_c1[22] ), .\nY_c1[23] (\nY_c1[23] ), 
            .\nY_c1[24] (\nY_c1[24] ), .\nY_c1[25] (\nY_c1[25] ), .\nY_c1[26] (\nY_c1[26] ), 
            .\nY1_c1[7] (\nY1_c1[7] ), .\nEY1_c1[9] (\nEY1_c1[9] ), .\nEY1_c1[10] (\nEY1_c1[10] ), 
            .\nEY1_c1[11] (\nEY1_c1[11] ), .\nEY1_c1[12] (\nEY1_c1[12] ), 
            .\nEY1_c1[13] (\nEY1_c1[13] ), .\nEY1_c1[14] (\nEY1_c1[14] ), 
            .\nEY1_c1[15] (\nEY1_c1[15] ), .\nEY1_c1[16] (\nEY1_c1[16] ), 
            .\nEY1_c1[17] (\nEY1_c1[17] ), .\nEY1_c1[0] (\nEY1_c1[0] ), 
            .\nEY1_c1[1] (\nEY1_c1[1] ), .\nEY1_c1[2] (\nEY1_c1[2] ), .\nEY1_c1[3] (\nEY1_c1[3] ), 
            .\nEY1_c1[4] (\nEY1_c1[4] ), .\nEY1_c1[5] (\nEY1_c1[5] ), .\nEY1_c1[6] (\nEY1_c1[6] ), 
            .\nEY1_c1[7] (\nEY1_c1[7] ), .\nEY1_c1[8] (\nEY1_c1[8] ), .clock(clock), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\nY_c1[10] (\nY_c1[10] ), 
            .\nY_c1[13] (\nY_c1[13] ), .\nY_c1[12] (\nY_c1[12] ), .\nEY1_c1[19] (\nEY1_c1[19] ), 
            .\nEY1_c1[20] (\nEY1_c1[20] ), .\nEY1_c1[21] (\nEY1_c1[21] ), 
            .\nEY1_c1[22] (\nEY1_c1[22] ), .\nEY1_c1[23] (\nEY1_c1[23] ), 
            .\nEY1_c1[24] (\nEY1_c1[24] ), .\nEY1_c1[18] (\nEY1_c1[18] ), 
            .\nY_c1[19] (\nY_c1[19] ), .\nY_c1[18] (\nY_c1[18] ), .\nY_c1[17] (\nY_c1[17] ), 
            .\nY_c1[16] (\nY_c1[16] ), .\nY_c1[15] (\nY_c1[15] ), .\nY_c1[14] (\nY_c1[14] ), 
            .\r0_1[13] (r0_1[13]), .\r0_1[11] (r0_1[11]), .\r0_1[12] (r0_1[12]), 
            .\r0_1[9] (r0_1[9]), .\r0_1[10] (r0_1[10]), .\r0_1[7] (r0_1[7]), 
            .\r0_1[8] (r0_1[8]), .\nY_c1[11] (\nY_c1[11] ), .\nY_c1[9] (\nY_c1[9] ), 
            .\buf_x[89] (\buf_x[89] ), .\s_1[0] (s_1[0]), .\buf_x[87] (\buf_x[87] ), 
            .\buf_x[88] (\buf_x[88] ), .\buf_x[85] (\buf_x[85] ), .\buf_x[86] (\buf_x[86] ), 
            .\buf_x[83] (\buf_x[83] ), .\buf_x[84] (\buf_x[84] ), .n70818(n70818), 
            .\buf_r[89] (\buf_r[89] ), .\buf_r[87] (\buf_r[87] ), .\buf_r[88] (\buf_r[88] ), 
            .\buf_r[85] (\buf_r[85] ), .\buf_r[86] (\buf_r[86] ), .\buf_r[83] (\buf_r[83] ), 
            .\buf_r[84] (\buf_r[84] ));
    
endmodule
//
// Verilog Description of module \mult_clk(8,6,false,false,1,3) 
//

module \mult_clk(8,6,false,false,1,3)  (\nY_c1[20] , \nY_c1[21] , \nY_c1[22] , 
            \nY_c1[23] , \nY_c1[24] , \nY_c1[25] , \nY_c1[26] , \nY1_c1[7] , 
            \nEY1_c1[9] , \nEY1_c1[10] , \nEY1_c1[11] , \nEY1_c1[12] , 
            \nEY1_c1[13] , \nEY1_c1[14] , \nEY1_c1[15] , \nEY1_c1[16] , 
            \nEY1_c1[17] , \nEY1_c1[0] , \nEY1_c1[1] , \nEY1_c1[2] , 
            \nEY1_c1[3] , \nEY1_c1[4] , \nEY1_c1[5] , \nEY1_c1[6] , 
            \nEY1_c1[7] , \nEY1_c1[8] , clock, GND_net, VCC_net, \nY_c1[10] , 
            \nY_c1[13] , \nY_c1[12] , \nEY1_c1[19] , \nEY1_c1[20] , 
            \nEY1_c1[21] , \nEY1_c1[22] , \nEY1_c1[23] , \nEY1_c1[24] , 
            \nEY1_c1[18] , \nY_c1[19] , \nY_c1[18] , \nY_c1[17] , \nY_c1[16] , 
            \nY_c1[15] , \nY_c1[14] , \r0_1[13] , \r0_1[11] , \r0_1[12] , 
            \r0_1[9] , \r0_1[10] , \r0_1[7] , \r0_1[8] , \nY_c1[11] , 
            \nY_c1[9] , \buf_x[89] , \s_1[0] , \buf_x[87] , \buf_x[88] , 
            \buf_x[85] , \buf_x[86] , \buf_x[83] , \buf_x[84] , n70818, 
            \buf_r[89] , \buf_r[87] , \buf_r[88] , \buf_r[85] , \buf_r[86] , 
            \buf_r[83] , \buf_r[84] );
    input \nY_c1[20] ;
    input \nY_c1[21] ;
    input \nY_c1[22] ;
    input \nY_c1[23] ;
    input \nY_c1[24] ;
    input \nY_c1[25] ;
    input \nY_c1[26] ;
    input \nY1_c1[7] ;
    output \nEY1_c1[9] ;
    output \nEY1_c1[10] ;
    output \nEY1_c1[11] ;
    output \nEY1_c1[12] ;
    output \nEY1_c1[13] ;
    output \nEY1_c1[14] ;
    output \nEY1_c1[15] ;
    output \nEY1_c1[16] ;
    output \nEY1_c1[17] ;
    output \nEY1_c1[0] ;
    output \nEY1_c1[1] ;
    output \nEY1_c1[2] ;
    output \nEY1_c1[3] ;
    output \nEY1_c1[4] ;
    output \nEY1_c1[5] ;
    output \nEY1_c1[6] ;
    output \nEY1_c1[7] ;
    output \nEY1_c1[8] ;
    input clock;
    input GND_net;
    input VCC_net;
    input \nY_c1[10] ;
    input \nY_c1[13] ;
    input \nY_c1[12] ;
    output \nEY1_c1[19] ;
    output \nEY1_c1[20] ;
    output \nEY1_c1[21] ;
    output \nEY1_c1[22] ;
    output \nEY1_c1[23] ;
    output \nEY1_c1[24] ;
    output \nEY1_c1[18] ;
    input \nY_c1[19] ;
    input \nY_c1[18] ;
    input \nY_c1[17] ;
    input \nY_c1[16] ;
    input \nY_c1[15] ;
    input \nY_c1[14] ;
    output \r0_1[13] ;
    output \r0_1[11] ;
    output \r0_1[12] ;
    output \r0_1[9] ;
    output \r0_1[10] ;
    output \r0_1[7] ;
    output \r0_1[8] ;
    input \nY_c1[11] ;
    input \nY_c1[9] ;
    output \buf_x[89] ;
    input \s_1[0] ;
    output \buf_x[87] ;
    output \buf_x[88] ;
    output \buf_x[85] ;
    output \buf_x[86] ;
    output \buf_x[83] ;
    output \buf_x[84] ;
    input n70818;
    input \buf_r[89] ;
    input \buf_r[87] ;
    input \buf_r[88] ;
    input \buf_r[85] ;
    input \buf_r[86] ;
    input \buf_r[83] ;
    input \buf_r[84] ;
    
    wire [166:0]buf_x;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(336[10:15])
    wire [166:0]buf_r;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(337[10:15])
    
    wire n70824, n70823, n61754, n61753, n61752, n61751, n62204, 
        n62203, n62202, n62201, n62200, n62199, n21368, n62198, 
        n62197, n21364, n62120, n62119, n62118, n62117, n62083, 
        n62082, n62081, n62080;
    
    PDPW8KC mux_5060 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\nY_c1[20] ), .ADR5(\nY_c1[21] ), 
            .ADR6(\nY_c1[22] ), .ADR7(\nY_c1[23] ), .ADR8(\nY_c1[24] ), 
            .ADR9(\nY_c1[25] ), .ADR10(\nY_c1[26] ), .ADR11(\nY1_c1[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(clock), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO0(\nEY1_c1[9] ), .DO1(\nEY1_c1[10] ), .DO2(\nEY1_c1[11] ), 
            .DO3(\nEY1_c1[12] ), .DO4(\nEY1_c1[13] ), .DO5(\nEY1_c1[14] ), 
            .DO6(\nEY1_c1[15] ), .DO7(\nEY1_c1[16] ), .DO8(\nEY1_c1[17] ), 
            .DO9(\nEY1_c1[0] ), .DO10(\nEY1_c1[1] ), .DO11(\nEY1_c1[2] ), 
            .DO12(\nEY1_c1[3] ), .DO13(\nEY1_c1[4] ), .DO14(\nEY1_c1[5] ), 
            .DO15(\nEY1_c1[6] ), .DO16(\nEY1_c1[7] ), .DO17(\nEY1_c1[8] ));
    defparam mux_5060.DATA_WIDTH_W = 18;
    defparam mux_5060.DATA_WIDTH_R = 18;
    defparam mux_5060.REGMODE = "NOREG";
    defparam mux_5060.CSDECODE_W = "0b000";
    defparam mux_5060.CSDECODE_R = "0b000";
    defparam mux_5060.GSR = "DISABLED";
    defparam mux_5060.RESETMODE = "ASYNC";
    defparam mux_5060.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_5060.INIT_DATA = "STATIC";
    defparam mux_5060.INITVAL_00 = "0x122113FF802E2101C9BB0B67B3A84C29F2919B0C09BF13A1D22ACAC1BC770D1313EAD33095A22CBF";
    defparam mux_5060.INITVAL_01 = "0x214B309D5A32B761BF02057F62F65019A080431A2F1801A53505E3431C771DFF90A8B5376A6249C6";
    defparam mux_5060.INITVAL_02 = "0x081DE2B0460E47C31E7B15E3D3A3BD1EEF403FDD296720F2AE3548B1BC030291129BAF113D839185";
    defparam mux_5060.INITVAL_03 = "0x0C4082925E066E12418E0225C209473F6481E9583E2731E1913E6AE1F1C2002C8219BB036932594B";
    defparam mux_5060.INITVAL_04 = "0x33B7A0A38C2123138765103202855D00E1319D3E332D70CED627137019F21C90137E5E13A022FBE8";
    defparam mux_5060.INITVAL_05 = "0x04EB5149E924C1F3554F0657217C8229A773BF4A0EAF621D72356B9096C31DD8932B0507F311DA05";
    defparam mux_5060.INITVAL_06 = "0x06AD50F227180EE217222B4BD359B7006070B9A817492236BC300223D0BA0A87E1876626D6D35A89";
    defparam mux_5060.INITVAL_07 = "0x003FF00FF5023DC03FAB0635A08EE20C23A0FD5B1403C18AD81DD242371B298B3301E7372AD3EAFF";
    defparam mux_5060.INITVAL_08 = "0x395D731E7D2AF972491B1EB0219542147D5102B00C5CC09122064A704056024240100B0040100000";
    defparam mux_5060.INITVAL_09 = "0x3A3FA2A0D81A6B50B5873CD472EDEA21768149B8084D23C8AC3153D26A7E1C86612EEB09E05015AC";
    defparam mux_5060.INITVAL_0A = "0x0BA81322931943900F68294171223C3B9CF25AC6105163B8B8275A213BCA00B272E3B11C55D0B023";
    defparam mux_5060.INITVAL_0B = "0x36E901383E30C1C0EA222D2450C47A2C0B80C6F52D7270F144315411431637AB81BC1D0073C25C0C";
    defparam mux_5060.INITVAL_0C = "0x05EE817FFA2ABE53E29E1241C270523C738128C0294E200B9318CC8318760AE9324F153F9F21AF1E";
    defparam mux_5060.INITVAL_0D = "0x034870A21D11B3F19FE322FFC2CB7F37261024960E2141AACE27EBB35DCD047FB13D3A23D7D348BB";
    defparam mux_5060.INITVAL_0E = "0x3A353351D930CAB2D3BC2A6FF2866A271EE2698226D1727CA32981A2BF6F2F2973318637C303D28A";
    defparam mux_5060.INITVAL_0F = "0x36AC824DED13E2803B6C345AD25CDD180EF0B1D73EF87339F32910F1F4CD165210E1FF06B5900124";
    defparam mux_5060.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5060.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    LUT4 i10019_1_lut_2_lut (.A(\nY_c1[10] ), .B(\nY_c1[13] ), .Z(buf_x[92])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i10019_1_lut_2_lut.init = 16'h9999;
    LUT4 i1_2_lut_rep_854 (.A(\nY_c1[10] ), .B(\nY_c1[13] ), .Z(n70824)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_854.init = 16'h6666;
    LUT4 i10023_1_lut_2_lut (.A(\nY_c1[12] ), .B(\nY_c1[13] ), .Z(buf_x[103])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i10023_1_lut_2_lut.init = 16'h9999;
    LUT4 i1_2_lut_rep_853 (.A(\nY_c1[12] ), .B(\nY_c1[13] ), .Z(n70823)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_853.init = 16'h6666;
    FD1S3AX buf_r_92__68_i1 (.D(buf_x[92]), .CK(clock), .Q(buf_r[92]));
    defparam buf_r_92__68_i1.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i1 (.D(buf_x[103]), .CK(clock), .Q(buf_x[138]));
    defparam buf_r_103__57_i1.GSR = "DISABLED";
    PDPW8KC mux_5061 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
            .DI8(GND_net), .DI9(GND_net), .DI10(GND_net), .DI11(GND_net), 
            .DI12(GND_net), .DI13(GND_net), .DI14(GND_net), .DI15(GND_net), 
            .DI16(GND_net), .DI17(GND_net), .ADW0(GND_net), .ADW1(GND_net), 
            .ADW2(GND_net), .ADW3(GND_net), .ADW4(GND_net), .ADW5(GND_net), 
            .ADW6(GND_net), .ADW7(GND_net), .ADW8(GND_net), .BE0(GND_net), 
            .BE1(GND_net), .CEW(VCC_net), .CLKW(GND_net), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(\nY_c1[20] ), .ADR5(\nY_c1[21] ), 
            .ADR6(\nY_c1[22] ), .ADR7(\nY_c1[23] ), .ADR8(\nY_c1[24] ), 
            .ADR9(\nY_c1[25] ), .ADR10(\nY_c1[26] ), .ADR11(\nY1_c1[7] ), 
            .ADR12(GND_net), .CER(VCC_net), .OCER(VCC_net), .CLKR(clock), 
            .CSR0(GND_net), .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), 
            .DO9(\nEY1_c1[19] ), .DO10(\nEY1_c1[20] ), .DO11(\nEY1_c1[21] ), 
            .DO12(\nEY1_c1[22] ), .DO13(\nEY1_c1[23] ), .DO14(\nEY1_c1[24] ), 
            .DO15(\nEY1_c1[18] ));
    defparam mux_5061.DATA_WIDTH_W = 18;
    defparam mux_5061.DATA_WIDTH_R = 18;
    defparam mux_5061.REGMODE = "NOREG";
    defparam mux_5061.CSDECODE_W = "0b000";
    defparam mux_5061.CSDECODE_R = "0b000";
    defparam mux_5061.GSR = "DISABLED";
    defparam mux_5061.RESETMODE = "ASYNC";
    defparam mux_5061.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_5061.INIT_DATA = "STATIC";
    defparam mux_5061.INITVAL_00 = "0x00064000630002300062000220002100060000200005F0005E0001E0005D0001D0001C0005B0001B";
    defparam mux_5061.INITVAL_01 = "0x0002F0006E0006D0002D0006C0006B0002B0006A0006900029000680006700027000660006500025";
    defparam mux_5061.INITVAL_02 = "0x0007A00079000390003800077000760003600075000740003400033000720003200031000700006F";
    defparam mux_5061.INITVAL_03 = "0x0004600045000050000400043000420004100001000000007F0007E0003E0007D0007C0003C0003B";
    defparam mux_5061.INITVAL_04 = "0x00013000520005100050000100000F0004E0004D0004C0000C0000B0004A00049000480000800007";
    defparam mux_5061.INITVAL_05 = "0x00021000200001F0001E0005D0005C0005B0005A0001A00019000180005700056000550001500014";
    defparam mux_5061.INITVAL_06 = "0x0006F0006E0006D0006C0006B0006A0002A000290002800027000260002500064000630006200061";
    defparam mux_5061.INITVAL_07 = "0x0003F0003E0003D0003C0003B0003A00039000380003700036000350003400033000320003100030";
    defparam mux_5061.INITVAL_08 = "0x0000F0000E0000D0000C0000B0000A00009000080000700006000050000400003000020000100000";
    defparam mux_5061.INITVAL_09 = "0x000600005F0005E0005D0001C0001B0001A000190001800056000550005400053000520005100050";
    defparam mux_5061.INITVAL_0A = "0x000730003200031000300006E0006D0002C0002B0002A00068000670006600065000240002300022";
    defparam mux_5061.INITVAL_0B = "0x0000700006000440004300002000010007F0007E0003D0003C0007A0007900038000370003600074";
    defparam mux_5061.INITVAL_0C = "0x0005C0001B00059000180001700055000140001300051000500000F0004D0004C0000B0004900048";
    defparam mux_5061.INITVAL_0D = "0x0003300071000300006E0002D0006B0002A000290006700026000640002300022000600001F0005D";
    defparam mux_5061.INITVAL_0E = "0x0004A000090004700006000440000300041000000007E0003D0007B0003A00078000370007500034";
    defparam mux_5061.INITVAL_0F = "0x0002400062000210005F0005D0001C0005A0001900017000550001400052000110004F0000E0004C";
    defparam mux_5061.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_5061.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    FD1S3AX buf_r_92__68_i2 (.D(buf_x[93]), .CK(clock), .Q(buf_r[93]));
    defparam buf_r_92__68_i2.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i3 (.D(buf_x[94]), .CK(clock), .Q(buf_r[94]));
    defparam buf_r_92__68_i3.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i4 (.D(buf_x[95]), .CK(clock), .Q(buf_r[95]));
    defparam buf_r_92__68_i4.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i5 (.D(buf_x[96]), .CK(clock), .Q(buf_r[96]));
    defparam buf_r_92__68_i5.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i6 (.D(buf_x[97]), .CK(clock), .Q(buf_r[97]));
    defparam buf_r_92__68_i6.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i7 (.D(buf_x[98]), .CK(clock), .Q(buf_r[98]));
    defparam buf_r_92__68_i7.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i8 (.D(buf_x[99]), .CK(clock), .Q(buf_r[99]));
    defparam buf_r_92__68_i8.GSR = "DISABLED";
    FD1S3AX buf_r_92__68_i9 (.D(buf_x[100]), .CK(clock), .Q(buf_r[100]));
    defparam buf_r_92__68_i9.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i2 (.D(buf_x[104]), .CK(clock), .Q(buf_x[139]));
    defparam buf_r_103__57_i2.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i3 (.D(buf_x[105]), .CK(clock), .Q(buf_x[140]));
    defparam buf_r_103__57_i3.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i4 (.D(buf_x[106]), .CK(clock), .Q(buf_x[141]));
    defparam buf_r_103__57_i4.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i5 (.D(buf_x[107]), .CK(clock), .Q(buf_x[142]));
    defparam buf_r_103__57_i5.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i6 (.D(buf_x[108]), .CK(clock), .Q(buf_x[143]));
    defparam buf_r_103__57_i6.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i7 (.D(buf_x[109]), .CK(clock), .Q(buf_x[144]));
    defparam buf_r_103__57_i7.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i8 (.D(buf_x[110]), .CK(clock), .Q(buf_x[145]));
    defparam buf_r_103__57_i8.GSR = "DISABLED";
    FD1S3AX buf_r_103__57_i9 (.D(buf_x[111]), .CK(clock), .Q(buf_x[146]));
    defparam buf_r_103__57_i9.GSR = "DISABLED";
    CCU2D add_4697_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61754), 
          .S0(buf_x[111]));
    defparam add_4697_cout.INIT0 = 16'h0000;
    defparam add_4697_cout.INIT1 = 16'h0000;
    defparam add_4697_cout.INJECT1_0 = "NO";
    defparam add_4697_cout.INJECT1_1 = "NO";
    CCU2D add_4697_7 (.A0(\nY_c1[19] ), .B0(n70823), .C0(\nY_c1[18] ), 
          .D0(GND_net), .A1(\nY_c1[19] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n61753), .COUT(n61754), .S0(buf_x[109]), 
          .S1(buf_x[110]));
    defparam add_4697_7.INIT0 = 16'hd2d2;
    defparam add_4697_7.INIT1 = 16'hfaaa;
    defparam add_4697_7.INJECT1_0 = "NO";
    defparam add_4697_7.INJECT1_1 = "NO";
    CCU2D add_4697_5 (.A0(\nY_c1[17] ), .B0(n70823), .C0(\nY_c1[16] ), 
          .D0(GND_net), .A1(\nY_c1[18] ), .B1(n70823), .C1(\nY_c1[17] ), 
          .D1(GND_net), .CIN(n61752), .COUT(n61753), .S0(buf_x[107]), 
          .S1(buf_x[108]));
    defparam add_4697_5.INIT0 = 16'hd2d2;
    defparam add_4697_5.INIT1 = 16'hd2d2;
    defparam add_4697_5.INJECT1_0 = "NO";
    defparam add_4697_5.INJECT1_1 = "NO";
    CCU2D add_4697_3 (.A0(\nY_c1[15] ), .B0(n70823), .C0(\nY_c1[14] ), 
          .D0(GND_net), .A1(\nY_c1[16] ), .B1(n70823), .C1(\nY_c1[15] ), 
          .D1(GND_net), .CIN(n61751), .COUT(n61752), .S0(buf_x[105]), 
          .S1(buf_x[106]));
    defparam add_4697_3.INIT0 = 16'hd2d2;
    defparam add_4697_3.INIT1 = 16'hd2d2;
    defparam add_4697_3.INJECT1_0 = "NO";
    defparam add_4697_3.INJECT1_1 = "NO";
    CCU2D add_4697_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\nY_c1[14] ), .B1(n70823), .C1(GND_net), .D1(GND_net), 
          .COUT(n61751), .S1(buf_x[104]));
    defparam add_4697_1.INIT0 = 16'hF000;
    defparam add_4697_1.INIT1 = 16'hdddd;
    defparam add_4697_1.INJECT1_0 = "NO";
    defparam add_4697_1.INJECT1_1 = "NO";
    CCU2D add_4623_10 (.A0(buf_x[136]), .B0(buf_x[146]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62204), .S0(\r0_1[13] ));
    defparam add_4623_10.INIT0 = 16'h5666;
    defparam add_4623_10.INIT1 = 16'h0000;
    defparam add_4623_10.INJECT1_0 = "NO";
    defparam add_4623_10.INJECT1_1 = "NO";
    CCU2D add_4623_8 (.A0(buf_x[135]), .B0(buf_x[144]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[136]), .B1(buf_x[145]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62203), .COUT(n62204), .S0(\r0_1[11] ), 
          .S1(\r0_1[12] ));
    defparam add_4623_8.INIT0 = 16'h5666;
    defparam add_4623_8.INIT1 = 16'h5666;
    defparam add_4623_8.INJECT1_0 = "NO";
    defparam add_4623_8.INJECT1_1 = "NO";
    CCU2D add_4623_6 (.A0(buf_x[133]), .B0(buf_x[142]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[134]), .B1(buf_x[143]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62202), .COUT(n62203), .S0(\r0_1[9] ), 
          .S1(\r0_1[10] ));
    defparam add_4623_6.INIT0 = 16'h5666;
    defparam add_4623_6.INIT1 = 16'h5666;
    defparam add_4623_6.INJECT1_0 = "NO";
    defparam add_4623_6.INJECT1_1 = "NO";
    CCU2D add_4623_4 (.A0(buf_x[131]), .B0(buf_x[140]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[132]), .B1(buf_x[141]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62201), .COUT(n62202), .S0(\r0_1[7] ), 
          .S1(\r0_1[8] ));
    defparam add_4623_4.INIT0 = 16'h5666;
    defparam add_4623_4.INIT1 = 16'h5666;
    defparam add_4623_4.INJECT1_0 = "NO";
    defparam add_4623_4.INJECT1_1 = "NO";
    CCU2D add_4623_2 (.A0(buf_x[129]), .B0(buf_x[138]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_x[130]), .B1(buf_x[139]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62201));
    defparam add_4623_2.INIT0 = 16'h7000;
    defparam add_4623_2.INIT1 = 16'h5666;
    defparam add_4623_2.INJECT1_0 = "NO";
    defparam add_4623_2.INJECT1_1 = "NO";
    CCU2D add_4621_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62200), 
          .S0(buf_x[100]));
    defparam add_4621_cout.INIT0 = 16'h0000;
    defparam add_4621_cout.INIT1 = 16'h0000;
    defparam add_4621_cout.INJECT1_0 = "NO";
    defparam add_4621_cout.INJECT1_1 = "NO";
    CCU2D add_4621_7 (.A0(\nY_c1[18] ), .B0(n21368), .C0(\nY_c1[19] ), 
          .D0(buf_x[92]), .A1(\nY_c1[19] ), .B1(n21368), .C1(GND_net), 
          .D1(GND_net), .CIN(n62199), .COUT(n62200), .S0(buf_x[98]), 
          .S1(buf_x[99]));
    defparam add_4621_7.INIT0 = 16'hd222;
    defparam add_4621_7.INIT1 = 16'hd222;
    defparam add_4621_7.INJECT1_0 = "NO";
    defparam add_4621_7.INJECT1_1 = "NO";
    CCU2D add_4621_5 (.A0(\nY_c1[16] ), .B0(n21368), .C0(\nY_c1[17] ), 
          .D0(buf_x[92]), .A1(\nY_c1[17] ), .B1(n21368), .C1(\nY_c1[18] ), 
          .D1(buf_x[92]), .CIN(n62198), .COUT(n62199), .S0(buf_x[96]), 
          .S1(buf_x[97]));
    defparam add_4621_5.INIT0 = 16'hd222;
    defparam add_4621_5.INIT1 = 16'hd222;
    defparam add_4621_5.INJECT1_0 = "NO";
    defparam add_4621_5.INJECT1_1 = "NO";
    CCU2D add_4621_3 (.A0(\nY_c1[14] ), .B0(n21368), .C0(\nY_c1[15] ), 
          .D0(buf_x[92]), .A1(\nY_c1[15] ), .B1(n21368), .C1(\nY_c1[16] ), 
          .D1(buf_x[92]), .CIN(n62197), .COUT(n62198), .S0(buf_x[94]), 
          .S1(buf_x[95]));
    defparam add_4621_3.INIT0 = 16'hd222;
    defparam add_4621_3.INIT1 = 16'hd222;
    defparam add_4621_3.INJECT1_0 = "NO";
    defparam add_4621_3.INJECT1_1 = "NO";
    CCU2D add_4621_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\nY_c1[14] ), .B1(n70824), .C1(\nY_c1[11] ), .D1(\nY_c1[13] ), 
          .COUT(n62197), .S1(buf_x[93]));
    defparam add_4621_1.INIT0 = 16'hF000;
    defparam add_4621_1.INIT1 = 16'hd22d;
    defparam add_4621_1.INJECT1_0 = "NO";
    defparam add_4621_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(\nY_c1[9] ), .B(\nY_c1[13] ), .Z(n21364)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_844 (.A(\nY_c1[11] ), .B(\nY_c1[13] ), .Z(n21368)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_844.init = 16'h6666;
    CCU2D add_4620_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62120), 
          .S0(\buf_x[89] ));
    defparam add_4620_cout.INIT0 = 16'h0000;
    defparam add_4620_cout.INIT1 = 16'h0000;
    defparam add_4620_cout.INJECT1_0 = "NO";
    defparam add_4620_cout.INJECT1_1 = "NO";
    CCU2D add_4620_7 (.A0(\nY_c1[18] ), .B0(n21364), .C0(\nY_c1[19] ), 
          .D0(\s_1[0] ), .A1(\nY_c1[19] ), .B1(n21364), .C1(GND_net), 
          .D1(GND_net), .CIN(n62119), .COUT(n62120), .S0(\buf_x[87] ), 
          .S1(\buf_x[88] ));
    defparam add_4620_7.INIT0 = 16'hd222;
    defparam add_4620_7.INIT1 = 16'hd222;
    defparam add_4620_7.INJECT1_0 = "NO";
    defparam add_4620_7.INJECT1_1 = "NO";
    CCU2D add_4620_5 (.A0(\nY_c1[16] ), .B0(n21364), .C0(\nY_c1[17] ), 
          .D0(\s_1[0] ), .A1(\nY_c1[17] ), .B1(n21364), .C1(\nY_c1[18] ), 
          .D1(\s_1[0] ), .CIN(n62118), .COUT(n62119), .S0(\buf_x[85] ), 
          .S1(\buf_x[86] ));
    defparam add_4620_5.INIT0 = 16'hd222;
    defparam add_4620_5.INIT1 = 16'hd222;
    defparam add_4620_5.INJECT1_0 = "NO";
    defparam add_4620_5.INJECT1_1 = "NO";
    CCU2D add_4620_3 (.A0(\nY_c1[14] ), .B0(n21364), .C0(\nY_c1[15] ), 
          .D0(\s_1[0] ), .A1(\nY_c1[15] ), .B1(n21364), .C1(\nY_c1[16] ), 
          .D1(\s_1[0] ), .CIN(n62117), .COUT(n62118), .S0(\buf_x[83] ), 
          .S1(\buf_x[84] ));
    defparam add_4620_3.INIT0 = 16'hd222;
    defparam add_4620_3.INIT1 = 16'hd222;
    defparam add_4620_3.INJECT1_0 = "NO";
    defparam add_4620_3.INJECT1_1 = "NO";
    CCU2D add_4620_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\nY_c1[14] ), .B1(n70818), .C1(\nY_c1[9] ), .D1(\nY_c1[13] ), 
          .COUT(n62117));
    defparam add_4620_1.INIT0 = 16'hF000;
    defparam add_4620_1.INIT1 = 16'hd22d;
    defparam add_4620_1.INJECT1_0 = "NO";
    defparam add_4620_1.INJECT1_1 = "NO";
    CCU2D add_4698_10 (.A0(buf_r[100]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62083), 
          .S0(buf_x[135]), .S1(buf_x[136]));
    defparam add_4698_10.INIT0 = 16'hfaaa;
    defparam add_4698_10.INIT1 = 16'h0000;
    defparam add_4698_10.INJECT1_0 = "NO";
    defparam add_4698_10.INJECT1_1 = "NO";
    CCU2D add_4698_8 (.A0(\buf_r[89] ), .B0(buf_r[98]), .C0(GND_net), 
          .D0(GND_net), .A1(buf_r[99]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62082), .COUT(n62083), .S0(buf_x[133]), 
          .S1(buf_x[134]));
    defparam add_4698_8.INIT0 = 16'h5666;
    defparam add_4698_8.INIT1 = 16'hfaaa;
    defparam add_4698_8.INJECT1_0 = "NO";
    defparam add_4698_8.INJECT1_1 = "NO";
    CCU2D add_4698_6 (.A0(\buf_r[87] ), .B0(buf_r[96]), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_r[88] ), .B1(buf_r[97]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62081), .COUT(n62082), .S0(buf_x[131]), 
          .S1(buf_x[132]));
    defparam add_4698_6.INIT0 = 16'h5666;
    defparam add_4698_6.INIT1 = 16'h5666;
    defparam add_4698_6.INJECT1_0 = "NO";
    defparam add_4698_6.INJECT1_1 = "NO";
    CCU2D add_4698_4 (.A0(\buf_r[85] ), .B0(buf_r[94]), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_r[86] ), .B1(buf_r[95]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62080), .COUT(n62081), .S0(buf_x[129]), 
          .S1(buf_x[130]));
    defparam add_4698_4.INIT0 = 16'h5666;
    defparam add_4698_4.INIT1 = 16'h5666;
    defparam add_4698_4.INJECT1_0 = "NO";
    defparam add_4698_4.INJECT1_1 = "NO";
    CCU2D add_4698_2 (.A0(\buf_r[83] ), .B0(buf_r[92]), .C0(GND_net), 
          .D0(GND_net), .A1(\buf_r[84] ), .B1(buf_r[93]), .C1(GND_net), 
          .D1(GND_net), .COUT(n62080));
    defparam add_4698_2.INIT0 = 16'h7000;
    defparam add_4698_2.INIT1 = 16'h5666;
    defparam add_4698_2.INJECT1_0 = "NO";
    defparam add_4698_2.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \fp_exp_exp_y1(23) 
//

module \fp_exp_exp_y1(23)  (\nX_c1[27] , \nKLog2_c1[34] , GND_net, \nY_c1[27] , 
            \nX_c1[25] , \nKLog2_c1[32] , \nX_c1[26] , \nKLog2_c1[33] , 
            \nY_c1[25] , \nY_c1[26] , \nX_c1[23] , \nKLog2_c1[30] , 
            \nX_c1[24] , \nKLog2_c1[31] , \nY_c1[23] , \nY_c1[24] , 
            \nX_c1[21] , \nKLog2_c1[28] , \nX_c1[22] , \nKLog2_c1[29] , 
            \nY_c1[21] , \nY_c1[22] , \nX_c1[19] , \nKLog2_c1[26] , 
            \nX_c1[20] , \nKLog2_c1[27] , \nY_c1[19] , \nY_c1[20] , 
            \nX_c1[17] , \nKLog2_c1[24] , \nX_c1[18] , \nKLog2_c1[25] , 
            \nY_c1[17] , \nY_c1[18] , \nX_c1[15] , \nKLog2_c1[22] , 
            \nX_c1[16] , \nKLog2_c1[23] , \nY_c1[15] , \nY_c1[16] , 
            \nX_c1[13] , \nKLog2_c1[20] , \nX_c1[14] , \nKLog2_c1[21] , 
            \nY_c1[13] , \nY_c1[14] , \nX_c1[11] , \nKLog2_c1[18] , 
            \nX_c1[12] , \nKLog2_c1[19] , \nY_c1[11] , \nY_c1[12] , 
            \nX_c1[9] , \nKLog2_c1[16] , \nX_c1[10] , \nKLog2_c1[17] , 
            \nY_c1[9] , \nY_c1[10] , \nX_c1[7] , \nKLog2_c1[14] , \nX_c1[8] , 
            \nKLog2_c1[15] , \nY_c1[7] , \nY_c1[8] , \nX_c1[5] , \nKLog2_c1[12] , 
            \nX_c1[6] , \nKLog2_c1[13] , \nY_c1[5] , \nY_c1[6] , \nX_c1[3] , 
            \nKLog2_c1[10] , \nX_c1[4] , \nKLog2_c1[11] , \nY_c1[3] , 
            \nY_c1[4] , \nX_c1[1] , \nKLog2_c1[8] , \nX_c1[2] , \nKLog2_c1[9] , 
            \nY_c1[1] , \nY_c1[2] , \nX_c1[0] , \nKLog2_c1[7] , \nY_c1[0] , 
            \nEY1_c1[25] , n62787);
    input \nX_c1[27] ;
    input \nKLog2_c1[34] ;
    input GND_net;
    output \nY_c1[27] ;
    input \nX_c1[25] ;
    input \nKLog2_c1[32] ;
    input \nX_c1[26] ;
    input \nKLog2_c1[33] ;
    output \nY_c1[25] ;
    output \nY_c1[26] ;
    input \nX_c1[23] ;
    input \nKLog2_c1[30] ;
    input \nX_c1[24] ;
    input \nKLog2_c1[31] ;
    output \nY_c1[23] ;
    output \nY_c1[24] ;
    input \nX_c1[21] ;
    input \nKLog2_c1[28] ;
    input \nX_c1[22] ;
    input \nKLog2_c1[29] ;
    output \nY_c1[21] ;
    output \nY_c1[22] ;
    input \nX_c1[19] ;
    input \nKLog2_c1[26] ;
    input \nX_c1[20] ;
    input \nKLog2_c1[27] ;
    output \nY_c1[19] ;
    output \nY_c1[20] ;
    input \nX_c1[17] ;
    input \nKLog2_c1[24] ;
    input \nX_c1[18] ;
    input \nKLog2_c1[25] ;
    output \nY_c1[17] ;
    output \nY_c1[18] ;
    input \nX_c1[15] ;
    input \nKLog2_c1[22] ;
    input \nX_c1[16] ;
    input \nKLog2_c1[23] ;
    output \nY_c1[15] ;
    output \nY_c1[16] ;
    input \nX_c1[13] ;
    input \nKLog2_c1[20] ;
    input \nX_c1[14] ;
    input \nKLog2_c1[21] ;
    output \nY_c1[13] ;
    output \nY_c1[14] ;
    input \nX_c1[11] ;
    input \nKLog2_c1[18] ;
    input \nX_c1[12] ;
    input \nKLog2_c1[19] ;
    output \nY_c1[11] ;
    output \nY_c1[12] ;
    input \nX_c1[9] ;
    input \nKLog2_c1[16] ;
    input \nX_c1[10] ;
    input \nKLog2_c1[17] ;
    output \nY_c1[9] ;
    output \nY_c1[10] ;
    input \nX_c1[7] ;
    input \nKLog2_c1[14] ;
    input \nX_c1[8] ;
    input \nKLog2_c1[15] ;
    output \nY_c1[7] ;
    output \nY_c1[8] ;
    input \nX_c1[5] ;
    input \nKLog2_c1[12] ;
    input \nX_c1[6] ;
    input \nKLog2_c1[13] ;
    output \nY_c1[5] ;
    output \nY_c1[6] ;
    input \nX_c1[3] ;
    input \nKLog2_c1[10] ;
    input \nX_c1[4] ;
    input \nKLog2_c1[11] ;
    output \nY_c1[3] ;
    output \nY_c1[4] ;
    input \nX_c1[1] ;
    input \nKLog2_c1[8] ;
    input \nX_c1[2] ;
    input \nKLog2_c1[9] ;
    output \nY_c1[1] ;
    output \nY_c1[2] ;
    input \nX_c1[0] ;
    input \nKLog2_c1[7] ;
    output \nY_c1[0] ;
    output \nEY1_c1[25] ;
    output n62787;
    
    
    fp_exp_exp_y1_23 \exp_y1_23.exp_y1  (.\nX_c1[27] (\nX_c1[27] ), .\nKLog2_c1[34] (\nKLog2_c1[34] ), 
            .GND_net(GND_net), .\nY_c1[27] (\nY_c1[27] ), .\nX_c1[25] (\nX_c1[25] ), 
            .\nKLog2_c1[32] (\nKLog2_c1[32] ), .\nX_c1[26] (\nX_c1[26] ), 
            .\nKLog2_c1[33] (\nKLog2_c1[33] ), .\nY_c1[25] (\nY_c1[25] ), 
            .\nY_c1[26] (\nY_c1[26] ), .\nX_c1[23] (\nX_c1[23] ), .\nKLog2_c1[30] (\nKLog2_c1[30] ), 
            .\nX_c1[24] (\nX_c1[24] ), .\nKLog2_c1[31] (\nKLog2_c1[31] ), 
            .\nY_c1[23] (\nY_c1[23] ), .\nY_c1[24] (\nY_c1[24] ), .\nX_c1[21] (\nX_c1[21] ), 
            .\nKLog2_c1[28] (\nKLog2_c1[28] ), .\nX_c1[22] (\nX_c1[22] ), 
            .\nKLog2_c1[29] (\nKLog2_c1[29] ), .\nY_c1[21] (\nY_c1[21] ), 
            .\nY_c1[22] (\nY_c1[22] ), .\nX_c1[19] (\nX_c1[19] ), .\nKLog2_c1[26] (\nKLog2_c1[26] ), 
            .\nX_c1[20] (\nX_c1[20] ), .\nKLog2_c1[27] (\nKLog2_c1[27] ), 
            .\nY_c1[19] (\nY_c1[19] ), .\nY_c1[20] (\nY_c1[20] ), .\nX_c1[17] (\nX_c1[17] ), 
            .\nKLog2_c1[24] (\nKLog2_c1[24] ), .\nX_c1[18] (\nX_c1[18] ), 
            .\nKLog2_c1[25] (\nKLog2_c1[25] ), .\nY_c1[17] (\nY_c1[17] ), 
            .\nY_c1[18] (\nY_c1[18] ), .\nX_c1[15] (\nX_c1[15] ), .\nKLog2_c1[22] (\nKLog2_c1[22] ), 
            .\nX_c1[16] (\nX_c1[16] ), .\nKLog2_c1[23] (\nKLog2_c1[23] ), 
            .\nY_c1[15] (\nY_c1[15] ), .\nY_c1[16] (\nY_c1[16] ), .\nX_c1[13] (\nX_c1[13] ), 
            .\nKLog2_c1[20] (\nKLog2_c1[20] ), .\nX_c1[14] (\nX_c1[14] ), 
            .\nKLog2_c1[21] (\nKLog2_c1[21] ), .\nY_c1[13] (\nY_c1[13] ), 
            .\nY_c1[14] (\nY_c1[14] ), .\nX_c1[11] (\nX_c1[11] ), .\nKLog2_c1[18] (\nKLog2_c1[18] ), 
            .\nX_c1[12] (\nX_c1[12] ), .\nKLog2_c1[19] (\nKLog2_c1[19] ), 
            .\nY_c1[11] (\nY_c1[11] ), .\nY_c1[12] (\nY_c1[12] ), .\nX_c1[9] (\nX_c1[9] ), 
            .\nKLog2_c1[16] (\nKLog2_c1[16] ), .\nX_c1[10] (\nX_c1[10] ), 
            .\nKLog2_c1[17] (\nKLog2_c1[17] ), .\nY_c1[9] (\nY_c1[9] ), 
            .\nY_c1[10] (\nY_c1[10] ), .\nX_c1[7] (\nX_c1[7] ), .\nKLog2_c1[14] (\nKLog2_c1[14] ), 
            .\nX_c1[8] (\nX_c1[8] ), .\nKLog2_c1[15] (\nKLog2_c1[15] ), 
            .\nY_c1[7] (\nY_c1[7] ), .\nY_c1[8] (\nY_c1[8] ), .\nX_c1[5] (\nX_c1[5] ), 
            .\nKLog2_c1[12] (\nKLog2_c1[12] ), .\nX_c1[6] (\nX_c1[6] ), 
            .\nKLog2_c1[13] (\nKLog2_c1[13] ), .\nY_c1[5] (\nY_c1[5] ), 
            .\nY_c1[6] (\nY_c1[6] ), .\nX_c1[3] (\nX_c1[3] ), .\nKLog2_c1[10] (\nKLog2_c1[10] ), 
            .\nX_c1[4] (\nX_c1[4] ), .\nKLog2_c1[11] (\nKLog2_c1[11] ), 
            .\nY_c1[3] (\nY_c1[3] ), .\nY_c1[4] (\nY_c1[4] ), .\nX_c1[1] (\nX_c1[1] ), 
            .\nKLog2_c1[8] (\nKLog2_c1[8] ), .\nX_c1[2] (\nX_c1[2] ), .\nKLog2_c1[9] (\nKLog2_c1[9] ), 
            .\nY_c1[1] (\nY_c1[1] ), .\nY_c1[2] (\nY_c1[2] ), .\nX_c1[0] (\nX_c1[0] ), 
            .\nKLog2_c1[7] (\nKLog2_c1[7] ), .\nY_c1[0] (\nY_c1[0] ), .\nEY1_c1[25] (\nEY1_c1[25] ), 
            .n62787(n62787));
    
endmodule
//
// Verilog Description of module fp_exp_exp_y1_23
//

module fp_exp_exp_y1_23 (\nX_c1[27] , \nKLog2_c1[34] , GND_net, \nY_c1[27] , 
            \nX_c1[25] , \nKLog2_c1[32] , \nX_c1[26] , \nKLog2_c1[33] , 
            \nY_c1[25] , \nY_c1[26] , \nX_c1[23] , \nKLog2_c1[30] , 
            \nX_c1[24] , \nKLog2_c1[31] , \nY_c1[23] , \nY_c1[24] , 
            \nX_c1[21] , \nKLog2_c1[28] , \nX_c1[22] , \nKLog2_c1[29] , 
            \nY_c1[21] , \nY_c1[22] , \nX_c1[19] , \nKLog2_c1[26] , 
            \nX_c1[20] , \nKLog2_c1[27] , \nY_c1[19] , \nY_c1[20] , 
            \nX_c1[17] , \nKLog2_c1[24] , \nX_c1[18] , \nKLog2_c1[25] , 
            \nY_c1[17] , \nY_c1[18] , \nX_c1[15] , \nKLog2_c1[22] , 
            \nX_c1[16] , \nKLog2_c1[23] , \nY_c1[15] , \nY_c1[16] , 
            \nX_c1[13] , \nKLog2_c1[20] , \nX_c1[14] , \nKLog2_c1[21] , 
            \nY_c1[13] , \nY_c1[14] , \nX_c1[11] , \nKLog2_c1[18] , 
            \nX_c1[12] , \nKLog2_c1[19] , \nY_c1[11] , \nY_c1[12] , 
            \nX_c1[9] , \nKLog2_c1[16] , \nX_c1[10] , \nKLog2_c1[17] , 
            \nY_c1[9] , \nY_c1[10] , \nX_c1[7] , \nKLog2_c1[14] , \nX_c1[8] , 
            \nKLog2_c1[15] , \nY_c1[7] , \nY_c1[8] , \nX_c1[5] , \nKLog2_c1[12] , 
            \nX_c1[6] , \nKLog2_c1[13] , \nY_c1[5] , \nY_c1[6] , \nX_c1[3] , 
            \nKLog2_c1[10] , \nX_c1[4] , \nKLog2_c1[11] , \nY_c1[3] , 
            \nY_c1[4] , \nX_c1[1] , \nKLog2_c1[8] , \nX_c1[2] , \nKLog2_c1[9] , 
            \nY_c1[1] , \nY_c1[2] , \nX_c1[0] , \nKLog2_c1[7] , \nY_c1[0] , 
            \nEY1_c1[25] , n62787);
    input \nX_c1[27] ;
    input \nKLog2_c1[34] ;
    input GND_net;
    output \nY_c1[27] ;
    input \nX_c1[25] ;
    input \nKLog2_c1[32] ;
    input \nX_c1[26] ;
    input \nKLog2_c1[33] ;
    output \nY_c1[25] ;
    output \nY_c1[26] ;
    input \nX_c1[23] ;
    input \nKLog2_c1[30] ;
    input \nX_c1[24] ;
    input \nKLog2_c1[31] ;
    output \nY_c1[23] ;
    output \nY_c1[24] ;
    input \nX_c1[21] ;
    input \nKLog2_c1[28] ;
    input \nX_c1[22] ;
    input \nKLog2_c1[29] ;
    output \nY_c1[21] ;
    output \nY_c1[22] ;
    input \nX_c1[19] ;
    input \nKLog2_c1[26] ;
    input \nX_c1[20] ;
    input \nKLog2_c1[27] ;
    output \nY_c1[19] ;
    output \nY_c1[20] ;
    input \nX_c1[17] ;
    input \nKLog2_c1[24] ;
    input \nX_c1[18] ;
    input \nKLog2_c1[25] ;
    output \nY_c1[17] ;
    output \nY_c1[18] ;
    input \nX_c1[15] ;
    input \nKLog2_c1[22] ;
    input \nX_c1[16] ;
    input \nKLog2_c1[23] ;
    output \nY_c1[15] ;
    output \nY_c1[16] ;
    input \nX_c1[13] ;
    input \nKLog2_c1[20] ;
    input \nX_c1[14] ;
    input \nKLog2_c1[21] ;
    output \nY_c1[13] ;
    output \nY_c1[14] ;
    input \nX_c1[11] ;
    input \nKLog2_c1[18] ;
    input \nX_c1[12] ;
    input \nKLog2_c1[19] ;
    output \nY_c1[11] ;
    output \nY_c1[12] ;
    input \nX_c1[9] ;
    input \nKLog2_c1[16] ;
    input \nX_c1[10] ;
    input \nKLog2_c1[17] ;
    output \nY_c1[9] ;
    output \nY_c1[10] ;
    input \nX_c1[7] ;
    input \nKLog2_c1[14] ;
    input \nX_c1[8] ;
    input \nKLog2_c1[15] ;
    output \nY_c1[7] ;
    output \nY_c1[8] ;
    input \nX_c1[5] ;
    input \nKLog2_c1[12] ;
    input \nX_c1[6] ;
    input \nKLog2_c1[13] ;
    output \nY_c1[5] ;
    output \nY_c1[6] ;
    input \nX_c1[3] ;
    input \nKLog2_c1[10] ;
    input \nX_c1[4] ;
    input \nKLog2_c1[11] ;
    output \nY_c1[3] ;
    output \nY_c1[4] ;
    input \nX_c1[1] ;
    input \nKLog2_c1[8] ;
    input \nX_c1[2] ;
    input \nKLog2_c1[9] ;
    output \nY_c1[1] ;
    output \nY_c1[2] ;
    input \nX_c1[0] ;
    input \nKLog2_c1[7] ;
    output \nY_c1[0] ;
    output \nEY1_c1[25] ;
    output n62787;
    
    
    wire n62563, n62562, n62561, n62560, n62559, n62558, n62557, 
        n62556, n62555, n62554, n62553, n62552, n62551, n62550, 
        n67566, n67564, n67565, n17, n62815;
    
    CCU2D sub_14_add_2_29 (.A0(\nX_c1[27] ), .B0(\nKLog2_c1[34] ), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62563), .S0(\nY_c1[27] ));
    defparam sub_14_add_2_29.INIT0 = 16'h5999;
    defparam sub_14_add_2_29.INIT1 = 16'h0000;
    defparam sub_14_add_2_29.INJECT1_0 = "NO";
    defparam sub_14_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_27 (.A0(\nX_c1[25] ), .B0(\nKLog2_c1[32] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[26] ), .B1(\nKLog2_c1[33] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62562), .COUT(n62563), .S0(\nY_c1[25] ), 
          .S1(\nY_c1[26] ));
    defparam sub_14_add_2_27.INIT0 = 16'h5999;
    defparam sub_14_add_2_27.INIT1 = 16'h5999;
    defparam sub_14_add_2_27.INJECT1_0 = "NO";
    defparam sub_14_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_25 (.A0(\nX_c1[23] ), .B0(\nKLog2_c1[30] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[24] ), .B1(\nKLog2_c1[31] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62561), .COUT(n62562), .S0(\nY_c1[23] ), 
          .S1(\nY_c1[24] ));
    defparam sub_14_add_2_25.INIT0 = 16'h5999;
    defparam sub_14_add_2_25.INIT1 = 16'h5999;
    defparam sub_14_add_2_25.INJECT1_0 = "NO";
    defparam sub_14_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_23 (.A0(\nX_c1[21] ), .B0(\nKLog2_c1[28] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[22] ), .B1(\nKLog2_c1[29] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62560), .COUT(n62561), .S0(\nY_c1[21] ), 
          .S1(\nY_c1[22] ));
    defparam sub_14_add_2_23.INIT0 = 16'h5999;
    defparam sub_14_add_2_23.INIT1 = 16'h5999;
    defparam sub_14_add_2_23.INJECT1_0 = "NO";
    defparam sub_14_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_21 (.A0(\nX_c1[19] ), .B0(\nKLog2_c1[26] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[20] ), .B1(\nKLog2_c1[27] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62559), .COUT(n62560), .S0(\nY_c1[19] ), 
          .S1(\nY_c1[20] ));
    defparam sub_14_add_2_21.INIT0 = 16'h5999;
    defparam sub_14_add_2_21.INIT1 = 16'h5999;
    defparam sub_14_add_2_21.INJECT1_0 = "NO";
    defparam sub_14_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_19 (.A0(\nX_c1[17] ), .B0(\nKLog2_c1[24] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[18] ), .B1(\nKLog2_c1[25] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62558), .COUT(n62559), .S0(\nY_c1[17] ), 
          .S1(\nY_c1[18] ));
    defparam sub_14_add_2_19.INIT0 = 16'h5999;
    defparam sub_14_add_2_19.INIT1 = 16'h5999;
    defparam sub_14_add_2_19.INJECT1_0 = "NO";
    defparam sub_14_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_17 (.A0(\nX_c1[15] ), .B0(\nKLog2_c1[22] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[16] ), .B1(\nKLog2_c1[23] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62557), .COUT(n62558), .S0(\nY_c1[15] ), 
          .S1(\nY_c1[16] ));
    defparam sub_14_add_2_17.INIT0 = 16'h5999;
    defparam sub_14_add_2_17.INIT1 = 16'h5999;
    defparam sub_14_add_2_17.INJECT1_0 = "NO";
    defparam sub_14_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_15 (.A0(\nX_c1[13] ), .B0(\nKLog2_c1[20] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[14] ), .B1(\nKLog2_c1[21] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62556), .COUT(n62557), .S0(\nY_c1[13] ), 
          .S1(\nY_c1[14] ));
    defparam sub_14_add_2_15.INIT0 = 16'h5999;
    defparam sub_14_add_2_15.INIT1 = 16'h5999;
    defparam sub_14_add_2_15.INJECT1_0 = "NO";
    defparam sub_14_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_13 (.A0(\nX_c1[11] ), .B0(\nKLog2_c1[18] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[12] ), .B1(\nKLog2_c1[19] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62555), .COUT(n62556), .S0(\nY_c1[11] ), 
          .S1(\nY_c1[12] ));
    defparam sub_14_add_2_13.INIT0 = 16'h5999;
    defparam sub_14_add_2_13.INIT1 = 16'h5999;
    defparam sub_14_add_2_13.INJECT1_0 = "NO";
    defparam sub_14_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_11 (.A0(\nX_c1[9] ), .B0(\nKLog2_c1[16] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[10] ), .B1(\nKLog2_c1[17] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62554), .COUT(n62555), .S0(\nY_c1[9] ), 
          .S1(\nY_c1[10] ));
    defparam sub_14_add_2_11.INIT0 = 16'h5999;
    defparam sub_14_add_2_11.INIT1 = 16'h5999;
    defparam sub_14_add_2_11.INJECT1_0 = "NO";
    defparam sub_14_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_9 (.A0(\nX_c1[7] ), .B0(\nKLog2_c1[14] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[8] ), .B1(\nKLog2_c1[15] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62553), .COUT(n62554), .S0(\nY_c1[7] ), 
          .S1(\nY_c1[8] ));
    defparam sub_14_add_2_9.INIT0 = 16'h5999;
    defparam sub_14_add_2_9.INIT1 = 16'h5999;
    defparam sub_14_add_2_9.INJECT1_0 = "NO";
    defparam sub_14_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_7 (.A0(\nX_c1[5] ), .B0(\nKLog2_c1[12] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[6] ), .B1(\nKLog2_c1[13] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62552), .COUT(n62553), .S0(\nY_c1[5] ), 
          .S1(\nY_c1[6] ));
    defparam sub_14_add_2_7.INIT0 = 16'h5999;
    defparam sub_14_add_2_7.INIT1 = 16'h5999;
    defparam sub_14_add_2_7.INJECT1_0 = "NO";
    defparam sub_14_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_5 (.A0(\nX_c1[3] ), .B0(\nKLog2_c1[10] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[4] ), .B1(\nKLog2_c1[11] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62551), .COUT(n62552), .S0(\nY_c1[3] ), 
          .S1(\nY_c1[4] ));
    defparam sub_14_add_2_5.INIT0 = 16'h5999;
    defparam sub_14_add_2_5.INIT1 = 16'h5999;
    defparam sub_14_add_2_5.INJECT1_0 = "NO";
    defparam sub_14_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_3 (.A0(\nX_c1[1] ), .B0(\nKLog2_c1[8] ), .C0(GND_net), 
          .D0(GND_net), .A1(\nX_c1[2] ), .B1(\nKLog2_c1[9] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62550), .COUT(n62551), .S0(\nY_c1[1] ), 
          .S1(\nY_c1[2] ));
    defparam sub_14_add_2_3.INIT0 = 16'h5999;
    defparam sub_14_add_2_3.INIT1 = 16'h5999;
    defparam sub_14_add_2_3.INJECT1_0 = "NO";
    defparam sub_14_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\nX_c1[0] ), .B1(\nKLog2_c1[7] ), .C1(GND_net), .D1(GND_net), 
          .COUT(n62550), .S1(\nY_c1[0] ));
    defparam sub_14_add_2_1.INIT0 = 16'h0000;
    defparam sub_14_add_2_1.INIT1 = 16'h5999;
    defparam sub_14_add_2_1.INJECT1_0 = "NO";
    defparam sub_14_add_2_1.INJECT1_1 = "NO";
    LUT4 i17921_3_lut (.A(\nY_c1[26] ), .B(n67566), .C(\nY_c1[25] ), .Z(\nEY1_c1[25] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17921_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut (.A(\nY_c1[23] ), .B(\nY_c1[26] ), .C(\nY_c1[24] ), 
         .D(\nY_c1[25] ), .Z(n62787)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'hc800;
    PFUMX i54655 (.BLUT(n67564), .ALUT(n67565), .C0(\nY_c1[23] ), .Z(n67566));
    LUT4 i1_2_lut (.A(\nY_c1[22] ), .B(\nY_c1[21] ), .Z(n17)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i54917_4_lut (.A(\nY_c1[26] ), .B(\nY_c1[24] ), .C(\nY_c1[27] ), 
         .D(n17), .Z(n67565)) /* synthesis lut_function=(A (C)+!A (B (C+(D)))) */ ;
    defparam i54917_4_lut.init = 16'he4e0;
    LUT4 i2_3_lut (.A(\nY_c1[21] ), .B(\nY_c1[20] ), .C(\nY_c1[22] ), 
         .Z(n62815)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i54653_4_lut (.A(\nY_c1[26] ), .B(\nY_c1[27] ), .C(\nY_c1[24] ), 
         .D(n62815), .Z(n67564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C (D)))) */ ;
    defparam i54653_4_lut.init = 16'hca8a;
    
endmodule
//
// Verilog Description of module \delay(22,1) 
//

module \delay(22,1)  (nZ0_d2, clock, \nZ0_d1[20] , \nZ0_d1[19] , \nZ0_d1[18] , 
            \nZ0_d1[17] , \nZ0_d1[16] , \nZ0_d1[15] , \nZ0_d1[14] , 
            \nZ0_d1[13] , \nZ0_d1[12] , \nZ0_d1[11] , \nZ0_d1[10] , 
            \nZ0_d1[9] , \nZ0_d1[8] , \nZ0_d1[7] , \nZ0_d1[6] , \nZ0_d1[5] , 
            \nZ0_d1[4] , \nZ0_d1[3] , \nZ0_d1[2] , \nZ0_d1[1] , \nEY2_d1[0] , 
            \nZ0_d1[21] , n23956, n23957, n23958, n23959, n23960, 
            n23961, n23962, n23963, n23964, n23965);
    output [21:0]nZ0_d2;
    input clock;
    input \nZ0_d1[20] ;
    input \nZ0_d1[19] ;
    input \nZ0_d1[18] ;
    input \nZ0_d1[17] ;
    input \nZ0_d1[16] ;
    input \nZ0_d1[15] ;
    input \nZ0_d1[14] ;
    input \nZ0_d1[13] ;
    input \nZ0_d1[12] ;
    input \nZ0_d1[11] ;
    input \nZ0_d1[10] ;
    input \nZ0_d1[9] ;
    input \nZ0_d1[8] ;
    input \nZ0_d1[7] ;
    input \nZ0_d1[6] ;
    input \nZ0_d1[5] ;
    input \nZ0_d1[4] ;
    input \nZ0_d1[3] ;
    input \nZ0_d1[2] ;
    input \nZ0_d1[1] ;
    input \nEY2_d1[0] ;
    input \nZ0_d1[21] ;
    output n23956;
    output n23957;
    output n23958;
    output n23959;
    output n23960;
    output n23961;
    output n23962;
    output n23963;
    output n23964;
    output n23965;
    
    
    FD1S3AX buf_42__27 (.D(\nZ0_d1[20] ), .CK(clock), .Q(nZ0_d2[20]));
    defparam buf_42__27.GSR = "DISABLED";
    FD1S3AX buf_41__28 (.D(\nZ0_d1[19] ), .CK(clock), .Q(nZ0_d2[19]));
    defparam buf_41__28.GSR = "DISABLED";
    FD1S3AX buf_40__29 (.D(\nZ0_d1[18] ), .CK(clock), .Q(nZ0_d2[18]));
    defparam buf_40__29.GSR = "DISABLED";
    FD1S3AX buf_39__30 (.D(\nZ0_d1[17] ), .CK(clock), .Q(nZ0_d2[17]));
    defparam buf_39__30.GSR = "DISABLED";
    FD1S3AX buf_38__31 (.D(\nZ0_d1[16] ), .CK(clock), .Q(nZ0_d2[16]));
    defparam buf_38__31.GSR = "DISABLED";
    FD1S3AX buf_37__32 (.D(\nZ0_d1[15] ), .CK(clock), .Q(nZ0_d2[15]));
    defparam buf_37__32.GSR = "DISABLED";
    FD1S3AX buf_36__33 (.D(\nZ0_d1[14] ), .CK(clock), .Q(nZ0_d2[14]));
    defparam buf_36__33.GSR = "DISABLED";
    FD1S3AX buf_35__34 (.D(\nZ0_d1[13] ), .CK(clock), .Q(nZ0_d2[13]));
    defparam buf_35__34.GSR = "DISABLED";
    FD1S3AX buf_34__35 (.D(\nZ0_d1[12] ), .CK(clock), .Q(nZ0_d2[12]));
    defparam buf_34__35.GSR = "DISABLED";
    FD1S3AX buf_33__36 (.D(\nZ0_d1[11] ), .CK(clock), .Q(nZ0_d2[11]));
    defparam buf_33__36.GSR = "DISABLED";
    FD1S3AX buf_32__37 (.D(\nZ0_d1[10] ), .CK(clock), .Q(nZ0_d2[10]));
    defparam buf_32__37.GSR = "DISABLED";
    FD1S3AX buf_31__38 (.D(\nZ0_d1[9] ), .CK(clock), .Q(nZ0_d2[9]));
    defparam buf_31__38.GSR = "DISABLED";
    FD1S3AX buf_30__39 (.D(\nZ0_d1[8] ), .CK(clock), .Q(nZ0_d2[8]));
    defparam buf_30__39.GSR = "DISABLED";
    FD1S3AX buf_29__40 (.D(\nZ0_d1[7] ), .CK(clock), .Q(nZ0_d2[7]));
    defparam buf_29__40.GSR = "DISABLED";
    FD1S3AX buf_28__41 (.D(\nZ0_d1[6] ), .CK(clock), .Q(nZ0_d2[6]));
    defparam buf_28__41.GSR = "DISABLED";
    FD1S3AX buf_27__42 (.D(\nZ0_d1[5] ), .CK(clock), .Q(nZ0_d2[5]));
    defparam buf_27__42.GSR = "DISABLED";
    FD1S3AX buf_26__43 (.D(\nZ0_d1[4] ), .CK(clock), .Q(nZ0_d2[4]));
    defparam buf_26__43.GSR = "DISABLED";
    FD1S3AX buf_25__44 (.D(\nZ0_d1[3] ), .CK(clock), .Q(nZ0_d2[3]));
    defparam buf_25__44.GSR = "DISABLED";
    FD1S3AX buf_24__45 (.D(\nZ0_d1[2] ), .CK(clock), .Q(nZ0_d2[2]));
    defparam buf_24__45.GSR = "DISABLED";
    FD1S3AX buf_23__46 (.D(\nZ0_d1[1] ), .CK(clock), .Q(nZ0_d2[1]));
    defparam buf_23__46.GSR = "DISABLED";
    FD1S3AX buf_22__47 (.D(\nEY2_d1[0] ), .CK(clock), .Q(nZ0_d2[0]));
    defparam buf_22__47.GSR = "DISABLED";
    FD1S3AX buf_43__26 (.D(\nZ0_d1[21] ), .CK(clock), .Q(nZ0_d2[21]));
    defparam buf_43__26.GSR = "DISABLED";
    LUT4 i12266_1_lut (.A(nZ0_d2[20]), .Z(n23956)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12266_1_lut.init = 16'h5555;
    LUT4 i12267_1_lut (.A(nZ0_d2[18]), .Z(n23957)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12267_1_lut.init = 16'h5555;
    LUT4 i12268_1_lut (.A(nZ0_d2[16]), .Z(n23958)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12268_1_lut.init = 16'h5555;
    LUT4 i12269_1_lut (.A(nZ0_d2[14]), .Z(n23959)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12269_1_lut.init = 16'h5555;
    LUT4 i12270_1_lut (.A(nZ0_d2[12]), .Z(n23960)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12270_1_lut.init = 16'h5555;
    LUT4 i12271_1_lut (.A(nZ0_d2[10]), .Z(n23961)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12271_1_lut.init = 16'h5555;
    LUT4 i12272_1_lut (.A(nZ0_d2[8]), .Z(n23962)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12272_1_lut.init = 16'h5555;
    LUT4 i12273_1_lut (.A(nZ0_d2[6]), .Z(n23963)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12273_1_lut.init = 16'h5555;
    LUT4 i12274_1_lut (.A(nZ0_d2[4]), .Z(n23964)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12274_1_lut.init = 16'h5555;
    LUT4 i12275_1_lut (.A(nZ0_d2[2]), .Z(n23965)) /* synthesis lut_function=(!(A)) */ ;
    defparam i12275_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \delay(36,2) 
//

module \delay(36,2)  (\buf[55] , \buf[53] , \buf[52] , \buf[51] , \buf[50] , 
            n65483, \r_0[10] , \buf[54] , \r_0[1] , \nY_d1[19] , clock, 
            \nY_d1[18] , \nY_d1[17] , \nY_d1[16] , \nY_d1[15] , \nY_d1[14] , 
            \nY_d1[13] , \nY_d1[12] , \nY_d1[11] , \nY_d1[10] , \nY_d1[9] , 
            \nY_d1[8] , \nY_d1[7] , \nY_d1[6] , \nY_d1[5] , \nY_d1[4] , 
            \nY_d1[3] , \nY_d1[2] , \nY_d1[1] , \nY_d1[0] , \nY_c1[19] , 
            \nY_c1[18] , \nY_c1[17] , \nY_c1[16] , \nY_c1[15] , \nY_c1[14] , 
            \nY_c1[13] , \nY_c1[12] , \nY_c1[11] , \nY_c1[10] , \nY_c1[9] , 
            \nY_c1[8] , \nY_c1[7] , \nY_c1[6] , \nY_c1[5] , \nY_c1[4] , 
            \nY_c1[3] , \nY_c1[2] , \nY_c1[1] , \nY_c1[0] , n62, \r_0[9] , 
            \r_0[4] , \r_0[0] , n70868, \r_0[3] , \r_0[5] , \r_0[2] );
    output \buf[55] ;
    output \buf[53] ;
    output \buf[52] ;
    output \buf[51] ;
    output \buf[50] ;
    output n65483;
    output \r_0[10] ;
    output \buf[54] ;
    output \r_0[1] ;
    output \nY_d1[19] ;
    input clock;
    output \nY_d1[18] ;
    output \nY_d1[17] ;
    output \nY_d1[16] ;
    output \nY_d1[15] ;
    output \nY_d1[14] ;
    output \nY_d1[13] ;
    output \nY_d1[12] ;
    output \nY_d1[11] ;
    output \nY_d1[10] ;
    output \nY_d1[9] ;
    output \nY_d1[8] ;
    output \nY_d1[7] ;
    output \nY_d1[6] ;
    output \nY_d1[5] ;
    output \nY_d1[4] ;
    output \nY_d1[3] ;
    output \nY_d1[2] ;
    output \nY_d1[1] ;
    output \nY_d1[0] ;
    input \nY_c1[19] ;
    input \nY_c1[18] ;
    input \nY_c1[17] ;
    input \nY_c1[16] ;
    input \nY_c1[15] ;
    input \nY_c1[14] ;
    input \nY_c1[13] ;
    input \nY_c1[12] ;
    input \nY_c1[11] ;
    input \nY_c1[10] ;
    input \nY_c1[9] ;
    input \nY_c1[8] ;
    input \nY_c1[7] ;
    input \nY_c1[6] ;
    input \nY_c1[5] ;
    input \nY_c1[4] ;
    input \nY_c1[3] ;
    input \nY_c1[2] ;
    input \nY_c1[1] ;
    input \nY_c1[0] ;
    output n62;
    output \r_0[9] ;
    output \r_0[4] ;
    output \r_0[0] ;
    output n70868;
    output \r_0[3] ;
    output \r_0[5] ;
    output \r_0[2] ;
    
    wire [107:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    
    wire n68700, n68701, n66778, n6, n67576, n67577, n68699, n70851, 
        n39616, n67621, n29970, n67567, n67568, n8, n29993, n67570, 
        n67571, n67573, n67574, n29978, n93, n71, n78, n65, 
        n97, n84, n68996, n68995, n68994, n68992, n68989, n68991, 
        n68990;
    
    LUT4 n68700_bdd_3_lut (.A(n68700), .B(\buf[55] ), .C(\buf[53] ), .Z(n68701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n68700_bdd_3_lut.init = 16'hcaca;
    LUT4 buf_53__bdd_4_lut_56039 (.A(\buf[52] ), .B(\buf[55] ), .C(\buf[51] ), 
         .D(\buf[50] ), .Z(n68700)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam buf_53__bdd_4_lut_56039.init = 16'hfbbb;
    PFUMX i24 (.BLUT(n66778), .ALUT(n6), .C0(\buf[53] ), .Z(n65483));
    PFUMX i54667 (.BLUT(n67576), .ALUT(n67577), .C0(\buf[52] ), .Z(\r_0[10] ));
    PFUMX i55269 (.BLUT(n68701), .ALUT(n68699), .C0(\buf[54] ), .Z(\r_0[1] ));
    FD1S3AX buf_91__92 (.D(\buf[55] ), .CK(clock), .Q(\nY_d1[19] ));
    defparam buf_91__92.GSR = "DISABLED";
    FD1S3AX buf_90__93 (.D(\buf[54] ), .CK(clock), .Q(\nY_d1[18] ));
    defparam buf_90__93.GSR = "DISABLED";
    FD1S3AX buf_89__94 (.D(\buf[53] ), .CK(clock), .Q(\nY_d1[17] ));
    defparam buf_89__94.GSR = "DISABLED";
    FD1S3AX buf_88__95 (.D(\buf[52] ), .CK(clock), .Q(\nY_d1[16] ));
    defparam buf_88__95.GSR = "DISABLED";
    FD1S3AX buf_87__96 (.D(\buf[51] ), .CK(clock), .Q(\nY_d1[15] ));
    defparam buf_87__96.GSR = "DISABLED";
    FD1S3AX buf_86__97 (.D(\buf[50] ), .CK(clock), .Q(\nY_d1[14] ));
    defparam buf_86__97.GSR = "DISABLED";
    FD1S3AX buf_85__98 (.D(\buf [49]), .CK(clock), .Q(\nY_d1[13] ));
    defparam buf_85__98.GSR = "DISABLED";
    FD1S3AX buf_84__99 (.D(\buf [48]), .CK(clock), .Q(\nY_d1[12] ));
    defparam buf_84__99.GSR = "DISABLED";
    FD1S3AX buf_83__100 (.D(\buf [47]), .CK(clock), .Q(\nY_d1[11] ));
    defparam buf_83__100.GSR = "DISABLED";
    FD1S3AX buf_82__101 (.D(\buf [46]), .CK(clock), .Q(\nY_d1[10] ));
    defparam buf_82__101.GSR = "DISABLED";
    FD1S3AX buf_81__102 (.D(\buf [45]), .CK(clock), .Q(\nY_d1[9] ));
    defparam buf_81__102.GSR = "DISABLED";
    FD1S3AX buf_80__103 (.D(\buf [44]), .CK(clock), .Q(\nY_d1[8] ));
    defparam buf_80__103.GSR = "DISABLED";
    FD1S3AX buf_79__104 (.D(\buf [43]), .CK(clock), .Q(\nY_d1[7] ));
    defparam buf_79__104.GSR = "DISABLED";
    FD1S3AX buf_78__105 (.D(\buf [42]), .CK(clock), .Q(\nY_d1[6] ));
    defparam buf_78__105.GSR = "DISABLED";
    FD1S3AX buf_77__106 (.D(\buf [41]), .CK(clock), .Q(\nY_d1[5] ));
    defparam buf_77__106.GSR = "DISABLED";
    FD1S3AX buf_76__107 (.D(\buf [40]), .CK(clock), .Q(\nY_d1[4] ));
    defparam buf_76__107.GSR = "DISABLED";
    FD1S3AX buf_75__108 (.D(\buf [39]), .CK(clock), .Q(\nY_d1[3] ));
    defparam buf_75__108.GSR = "DISABLED";
    FD1S3AX buf_74__109 (.D(\buf [38]), .CK(clock), .Q(\nY_d1[2] ));
    defparam buf_74__109.GSR = "DISABLED";
    FD1S3AX buf_73__110 (.D(\buf [37]), .CK(clock), .Q(\nY_d1[1] ));
    defparam buf_73__110.GSR = "DISABLED";
    FD1S3AX buf_72__111 (.D(\buf [36]), .CK(clock), .Q(\nY_d1[0] ));
    defparam buf_72__111.GSR = "DISABLED";
    FD1S3AX buf_55__128 (.D(\nY_c1[19] ), .CK(clock), .Q(\buf[55] ));
    defparam buf_55__128.GSR = "DISABLED";
    FD1S3AX buf_54__129 (.D(\nY_c1[18] ), .CK(clock), .Q(\buf[54] ));
    defparam buf_54__129.GSR = "DISABLED";
    FD1S3AX buf_53__130 (.D(\nY_c1[17] ), .CK(clock), .Q(\buf[53] ));
    defparam buf_53__130.GSR = "DISABLED";
    FD1S3AX buf_52__131 (.D(\nY_c1[16] ), .CK(clock), .Q(\buf[52] ));
    defparam buf_52__131.GSR = "DISABLED";
    FD1S3AX buf_51__132 (.D(\nY_c1[15] ), .CK(clock), .Q(\buf[51] ));
    defparam buf_51__132.GSR = "DISABLED";
    FD1S3AX buf_50__133 (.D(\nY_c1[14] ), .CK(clock), .Q(\buf[50] ));
    defparam buf_50__133.GSR = "DISABLED";
    FD1S3AX buf_49__134 (.D(\nY_c1[13] ), .CK(clock), .Q(\buf [49]));
    defparam buf_49__134.GSR = "DISABLED";
    FD1S3AX buf_48__135 (.D(\nY_c1[12] ), .CK(clock), .Q(\buf [48]));
    defparam buf_48__135.GSR = "DISABLED";
    FD1S3AX buf_47__136 (.D(\nY_c1[11] ), .CK(clock), .Q(\buf [47]));
    defparam buf_47__136.GSR = "DISABLED";
    FD1S3AX buf_46__137 (.D(\nY_c1[10] ), .CK(clock), .Q(\buf [46]));
    defparam buf_46__137.GSR = "DISABLED";
    FD1S3AX buf_45__138 (.D(\nY_c1[9] ), .CK(clock), .Q(\buf [45]));
    defparam buf_45__138.GSR = "DISABLED";
    FD1S3AX buf_44__139 (.D(\nY_c1[8] ), .CK(clock), .Q(\buf [44]));
    defparam buf_44__139.GSR = "DISABLED";
    FD1S3AX buf_43__140 (.D(\nY_c1[7] ), .CK(clock), .Q(\buf [43]));
    defparam buf_43__140.GSR = "DISABLED";
    FD1S3AX buf_42__141 (.D(\nY_c1[6] ), .CK(clock), .Q(\buf [42]));
    defparam buf_42__141.GSR = "DISABLED";
    FD1S3AX buf_41__142 (.D(\nY_c1[5] ), .CK(clock), .Q(\buf [41]));
    defparam buf_41__142.GSR = "DISABLED";
    FD1S3AX buf_40__143 (.D(\nY_c1[4] ), .CK(clock), .Q(\buf [40]));
    defparam buf_40__143.GSR = "DISABLED";
    FD1S3AX buf_39__144 (.D(\nY_c1[3] ), .CK(clock), .Q(\buf [39]));
    defparam buf_39__144.GSR = "DISABLED";
    FD1S3AX buf_38__145 (.D(\nY_c1[2] ), .CK(clock), .Q(\buf [38]));
    defparam buf_38__145.GSR = "DISABLED";
    FD1S3AX buf_37__146 (.D(\nY_c1[1] ), .CK(clock), .Q(\buf [37]));
    defparam buf_37__146.GSR = "DISABLED";
    FD1S3AX buf_36__147 (.D(\nY_c1[0] ), .CK(clock), .Q(\buf [36]));
    defparam buf_36__147.GSR = "DISABLED";
    LUT4 buf_54__bdd_2_lut (.A(\buf[53] ), .B(\buf[55] ), .Z(n68699)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam buf_54__bdd_2_lut.init = 16'h4444;
    LUT4 i124_4_lut (.A(n70851), .B(\buf[54] ), .C(\buf[52] ), .D(\buf[53] ), 
         .Z(n62)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i124_4_lut.init = 16'heccc;
    LUT4 i28024_2_lut (.A(\buf[54] ), .B(\buf[53] ), .Z(n39616)) /* synthesis lut_function=(A (B)) */ ;
    defparam i28024_2_lut.init = 16'h8888;
    LUT4 i55004_2_lut (.A(\buf[55] ), .B(\buf[54] ), .Z(n67621)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i55004_2_lut.init = 16'h6666;
    LUT4 i54665_4_lut (.A(\buf[51] ), .B(n67621), .C(\buf[53] ), .D(n29970), 
         .Z(n67576)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i54665_4_lut.init = 16'hcac0;
    L6MUX21 i54658 (.D0(n67567), .D1(n67568), .SD(\buf[52] ), .Z(\r_0[9] ));
    PFUMX i54657 (.BLUT(n8), .ALUT(n29993), .C0(\buf[53] ), .Z(n67568));
    PFUMX i54661 (.BLUT(n67570), .ALUT(n67571), .C0(\buf[52] ), .Z(\r_0[4] ));
    PFUMX i54664 (.BLUT(n67573), .ALUT(n67574), .C0(\buf[52] ), .Z(\r_0[0] ));
    PFUMX i54666 (.BLUT(n29978), .ALUT(n93), .C0(\buf[53] ), .Z(n67577));
    PFUMX i54656 (.BLUT(n71), .ALUT(n78), .C0(\buf[53] ), .Z(n67567));
    LUT4 i55046_3_lut_4_lut (.A(\buf[50] ), .B(\buf[55] ), .C(\buf[51] ), 
         .D(\buf[54] ), .Z(n8)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i55046_3_lut_4_lut.init = 16'h5b4c;
    LUT4 i1_3_lut_4_lut (.A(\buf[50] ), .B(\buf[55] ), .C(\buf[54] ), 
         .D(\buf[51] ), .Z(n93)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i18352_3_lut_4_lut_4_lut (.A(\buf[50] ), .B(\buf[55] ), .C(\buf[51] ), 
         .D(\buf[54] ), .Z(n29993)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i18352_3_lut_4_lut_4_lut.init = 16'hf304;
    LUT4 i54662_4_lut_4_lut (.A(\buf[55] ), .B(n65), .C(\buf[53] ), .D(\buf[54] ), 
         .Z(n67573)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;
    defparam i54662_4_lut_4_lut.init = 16'h5f5c;
    LUT4 i6_1_lut_rep_898 (.A(\buf[55] ), .Z(n70868)) /* synthesis lut_function=(!(A)) */ ;
    defparam i6_1_lut_rep_898.init = 16'h5555;
    LUT4 i1_2_lut_3_lut (.A(\buf[54] ), .B(\buf[55] ), .C(\buf[50] ), 
         .Z(n97)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i1_2_lut_3_lut_adj_840 (.A(\buf[54] ), .B(\buf[55] ), .C(\buf[50] ), 
         .Z(n84)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_840.init = 16'hf8f8;
    LUT4 n68997_bdd_3_lut_4_lut (.A(\buf[52] ), .B(\buf[51] ), .C(\buf[54] ), 
         .D(n68996), .Z(\r_0[3] )) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam n68997_bdd_3_lut_4_lut.init = 16'hf606;
    PFUMX i55360 (.BLUT(n68995), .ALUT(n68994), .C0(\buf[53] ), .Z(n68996));
    LUT4 buf_52__bdd_2_lut_55362 (.A(\buf[52] ), .B(\buf[51] ), .Z(n68995)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam buf_52__bdd_2_lut_55362.init = 16'h6666;
    LUT4 buf_52__bdd_4_lut_55885 (.A(\buf[52] ), .B(\buf[50] ), .C(\buf[51] ), 
         .D(\buf[55] ), .Z(n68994)) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam buf_52__bdd_4_lut_55885.init = 16'h665a;
    LUT4 n68992_bdd_3_lut (.A(n68992), .B(n68989), .C(\buf[50] ), .Z(\r_0[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n68992_bdd_3_lut.init = 16'hcaca;
    PFUMX i55357 (.BLUT(n68991), .ALUT(n68990), .C0(\buf[51] ), .Z(n68992));
    LUT4 buf_55__bdd_2_lut_55895 (.A(\buf[54] ), .B(\buf[52] ), .Z(n68991)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam buf_55__bdd_2_lut_55895.init = 16'h6666;
    LUT4 buf_50__bdd_4_lut_56043 (.A(\buf[54] ), .B(\buf[52] ), .C(\buf[53] ), 
         .D(\buf[51] ), .Z(n68989)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam buf_50__bdd_4_lut_56043.init = 16'h6656;
    LUT4 buf_55__bdd_4_lut_56042 (.A(\buf[55] ), .B(\buf[54] ), .C(\buf[52] ), 
         .D(\buf[53] ), .Z(n68990)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A (B (C (D))+!B !(C (D))))) */ ;
    defparam buf_55__bdd_4_lut_56042.init = 16'h34cc;
    LUT4 i1_2_lut (.A(\buf[51] ), .B(\buf[55] ), .Z(n78)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_841 (.A(\buf[51] ), .B(\buf[50] ), .C(\buf[55] ), 
         .Z(n65)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_841.init = 16'h7070;
    LUT4 i54659_4_lut_4_lut (.A(\buf[51] ), .B(\buf[50] ), .C(n84), .D(\buf[53] ), 
         .Z(n67570)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A !(D))) */ ;
    defparam i54659_4_lut_4_lut.init = 16'h5f88;
    LUT4 i53875_3_lut_4_lut (.A(\buf[51] ), .B(\buf[50] ), .C(\buf[52] ), 
         .D(\buf[54] ), .Z(n66778)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i53875_3_lut_4_lut.init = 16'h80ff;
    LUT4 i54660_4_lut_4_lut (.A(\buf[51] ), .B(\buf[50] ), .C(n97), .D(\buf[53] ), 
         .Z(n67571)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B (C (D))))) */ ;
    defparam i54660_4_lut_4_lut.init = 16'h50ee;
    LUT4 i55070_3_lut_4_lut (.A(\buf[51] ), .B(\buf[50] ), .C(\buf[54] ), 
         .D(\buf[52] ), .Z(n6)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i55070_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i1_2_lut_rep_881 (.A(\buf[51] ), .B(\buf[50] ), .Z(n70851)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_881.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_842 (.A(\buf[50] ), .B(\buf[55] ), .C(\buf[54] ), 
         .D(\buf[51] ), .Z(n71)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i1_3_lut_4_lut_adj_842.init = 16'h70f0;
    LUT4 i1_2_lut_3_lut_adj_843 (.A(\buf[50] ), .B(\buf[55] ), .C(\buf[54] ), 
         .Z(n29970)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_843.init = 16'h8080;
    LUT4 i32_4_lut_4_lut (.A(\buf[55] ), .B(\buf[50] ), .C(n39616), .D(\buf[51] ), 
         .Z(\r_0[2] )) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B !(D))) */ ;
    defparam i32_4_lut_4_lut.init = 16'h936c;
    LUT4 i54663_4_lut (.A(\buf[54] ), .B(\buf[55] ), .C(\buf[53] ), .D(n70851), 
         .Z(n67574)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(B+!(C))) */ ;
    defparam i54663_4_lut.init = 16'hba3a;
    LUT4 i18337_3_lut_4_lut_4_lut (.A(\buf[54] ), .B(\buf[55] ), .C(\buf[51] ), 
         .D(\buf[50] ), .Z(n29978)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (C (D))))) */ ;
    defparam i18337_3_lut_4_lut_4_lut.init = 16'h6888;
    
endmodule
//
// Verilog Description of module \delay(36,4) 
//

module \delay(36,4)  (\nX_c1[27] , clock, \nX_c1[26] , \nX_c1[25] , 
            \nX_c1[24] , \nX_c1[23] , \nX_c1[22] , \nX_c1[21] , \nX_c1[20] , 
            \nX_c1[19] , \nX_c1[18] , \nX_c1[17] , \nX_c1[16] , \nX_c1[15] , 
            \nX_c1[14] , \nX_c1[13] , \nX_c1[12] , \nX_c1[11] , \nX_c1[10] , 
            \nX_c1[9] , \nX_c1[8] , \nX_c1[7] , \nX_c1[6] , \nX_c1[5] , 
            \nX_c1[4] , \nX_c1[3] , \nX_c1[2] , \nX_c1[1] , \nX_c1[0] , 
            \buf_x[437] , \buf_x[436] , \buf_x[435] , \buf_x[434] , 
            \nX_a1[23] , \nX_a1[22] , \nX_a1[21] , \nX_a1[20] , \nX_a1[19] , 
            \nX_a1[18] , \nX_a1[17] , \nX_a1[16] , \nX_a1[15] , \nX_a1[14] , 
            \nX_a1[13] , \nX_a1[12] , \nX_a1[11] , \nX_a1[10] , \nX_a1[9] , 
            \nX_a1[8] , \nX_a1[7] , \nX_a1[6] , \nX_a1[5] , \nX_a1[4] , 
            \nX_a1[3] , \nX_a1[2] , \nX_a1[1] , \nX_a1[0] );
    output \nX_c1[27] ;
    input clock;
    output \nX_c1[26] ;
    output \nX_c1[25] ;
    output \nX_c1[24] ;
    output \nX_c1[23] ;
    output \nX_c1[22] ;
    output \nX_c1[21] ;
    output \nX_c1[20] ;
    output \nX_c1[19] ;
    output \nX_c1[18] ;
    output \nX_c1[17] ;
    output \nX_c1[16] ;
    output \nX_c1[15] ;
    output \nX_c1[14] ;
    output \nX_c1[13] ;
    output \nX_c1[12] ;
    output \nX_c1[11] ;
    output \nX_c1[10] ;
    output \nX_c1[9] ;
    output \nX_c1[8] ;
    output \nX_c1[7] ;
    output \nX_c1[6] ;
    output \nX_c1[5] ;
    output \nX_c1[4] ;
    output \nX_c1[3] ;
    output \nX_c1[2] ;
    output \nX_c1[1] ;
    output \nX_c1[0] ;
    input \buf_x[437] ;
    input \buf_x[436] ;
    input \buf_x[435] ;
    input \buf_x[434] ;
    input \nX_a1[23] ;
    input \nX_a1[22] ;
    input \nX_a1[21] ;
    input \nX_a1[20] ;
    input \nX_a1[19] ;
    input \nX_a1[18] ;
    input \nX_a1[17] ;
    input \nX_a1[16] ;
    input \nX_a1[15] ;
    input \nX_a1[14] ;
    input \nX_a1[13] ;
    input \nX_a1[12] ;
    input \nX_a1[11] ;
    input \nX_a1[10] ;
    input \nX_a1[9] ;
    input \nX_a1[8] ;
    input \nX_a1[7] ;
    input \nX_a1[6] ;
    input \nX_a1[5] ;
    input \nX_a1[4] ;
    input \nX_a1[3] ;
    input \nX_a1[2] ;
    input \nX_a1[1] ;
    input \nX_a1[0] ;
    
    wire [179:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    
    FD1S3AX buf_171__156 (.D(\buf [135]), .CK(clock), .Q(\nX_c1[27] ));
    defparam buf_171__156.GSR = "DISABLED";
    FD1S3AX buf_170__157 (.D(\buf [134]), .CK(clock), .Q(\nX_c1[26] ));
    defparam buf_170__157.GSR = "DISABLED";
    FD1S3AX buf_169__158 (.D(\buf [133]), .CK(clock), .Q(\nX_c1[25] ));
    defparam buf_169__158.GSR = "DISABLED";
    FD1S3AX buf_168__159 (.D(\buf [132]), .CK(clock), .Q(\nX_c1[24] ));
    defparam buf_168__159.GSR = "DISABLED";
    FD1S3AX buf_167__160 (.D(\buf [131]), .CK(clock), .Q(\nX_c1[23] ));
    defparam buf_167__160.GSR = "DISABLED";
    FD1S3AX buf_166__161 (.D(\buf [130]), .CK(clock), .Q(\nX_c1[22] ));
    defparam buf_166__161.GSR = "DISABLED";
    FD1S3AX buf_165__162 (.D(\buf [129]), .CK(clock), .Q(\nX_c1[21] ));
    defparam buf_165__162.GSR = "DISABLED";
    FD1S3AX buf_164__163 (.D(\buf [128]), .CK(clock), .Q(\nX_c1[20] ));
    defparam buf_164__163.GSR = "DISABLED";
    FD1S3AX buf_163__164 (.D(\buf [127]), .CK(clock), .Q(\nX_c1[19] ));
    defparam buf_163__164.GSR = "DISABLED";
    FD1S3AX buf_162__165 (.D(\buf [126]), .CK(clock), .Q(\nX_c1[18] ));
    defparam buf_162__165.GSR = "DISABLED";
    FD1S3AX buf_161__166 (.D(\buf [125]), .CK(clock), .Q(\nX_c1[17] ));
    defparam buf_161__166.GSR = "DISABLED";
    FD1S3AX buf_160__167 (.D(\buf [124]), .CK(clock), .Q(\nX_c1[16] ));
    defparam buf_160__167.GSR = "DISABLED";
    FD1S3AX buf_159__168 (.D(\buf [123]), .CK(clock), .Q(\nX_c1[15] ));
    defparam buf_159__168.GSR = "DISABLED";
    FD1S3AX buf_158__169 (.D(\buf [122]), .CK(clock), .Q(\nX_c1[14] ));
    defparam buf_158__169.GSR = "DISABLED";
    FD1S3AX buf_157__170 (.D(\buf [121]), .CK(clock), .Q(\nX_c1[13] ));
    defparam buf_157__170.GSR = "DISABLED";
    FD1S3AX buf_156__171 (.D(\buf [120]), .CK(clock), .Q(\nX_c1[12] ));
    defparam buf_156__171.GSR = "DISABLED";
    FD1S3AX buf_155__172 (.D(\buf [119]), .CK(clock), .Q(\nX_c1[11] ));
    defparam buf_155__172.GSR = "DISABLED";
    FD1S3AX buf_154__173 (.D(\buf [118]), .CK(clock), .Q(\nX_c1[10] ));
    defparam buf_154__173.GSR = "DISABLED";
    FD1S3AX buf_153__174 (.D(\buf [117]), .CK(clock), .Q(\nX_c1[9] ));
    defparam buf_153__174.GSR = "DISABLED";
    FD1S3AX buf_152__175 (.D(\buf [116]), .CK(clock), .Q(\nX_c1[8] ));
    defparam buf_152__175.GSR = "DISABLED";
    FD1S3AX buf_151__176 (.D(\buf [115]), .CK(clock), .Q(\nX_c1[7] ));
    defparam buf_151__176.GSR = "DISABLED";
    FD1S3AX buf_150__177 (.D(\buf [114]), .CK(clock), .Q(\nX_c1[6] ));
    defparam buf_150__177.GSR = "DISABLED";
    FD1S3AX buf_149__178 (.D(\buf [113]), .CK(clock), .Q(\nX_c1[5] ));
    defparam buf_149__178.GSR = "DISABLED";
    FD1S3AX buf_148__179 (.D(\buf [112]), .CK(clock), .Q(\nX_c1[4] ));
    defparam buf_148__179.GSR = "DISABLED";
    FD1S3AX buf_147__180 (.D(\buf [111]), .CK(clock), .Q(\nX_c1[3] ));
    defparam buf_147__180.GSR = "DISABLED";
    FD1S3AX buf_146__181 (.D(\buf [110]), .CK(clock), .Q(\nX_c1[2] ));
    defparam buf_146__181.GSR = "DISABLED";
    FD1S3AX buf_145__182 (.D(\buf [109]), .CK(clock), .Q(\nX_c1[1] ));
    defparam buf_145__182.GSR = "DISABLED";
    FD1S3AX buf_144__183 (.D(\buf [108]), .CK(clock), .Q(\nX_c1[0] ));
    defparam buf_144__183.GSR = "DISABLED";
    FD1S3AX buf_135__192 (.D(\buf [99]), .CK(clock), .Q(\buf [135]));
    defparam buf_135__192.GSR = "DISABLED";
    FD1S3AX buf_134__193 (.D(\buf [98]), .CK(clock), .Q(\buf [134]));
    defparam buf_134__193.GSR = "DISABLED";
    FD1S3AX buf_133__194 (.D(\buf [97]), .CK(clock), .Q(\buf [133]));
    defparam buf_133__194.GSR = "DISABLED";
    FD1S3AX buf_132__195 (.D(\buf [96]), .CK(clock), .Q(\buf [132]));
    defparam buf_132__195.GSR = "DISABLED";
    FD1S3AX buf_131__196 (.D(\buf [95]), .CK(clock), .Q(\buf [131]));
    defparam buf_131__196.GSR = "DISABLED";
    FD1S3AX buf_130__197 (.D(\buf [94]), .CK(clock), .Q(\buf [130]));
    defparam buf_130__197.GSR = "DISABLED";
    FD1S3AX buf_129__198 (.D(\buf [93]), .CK(clock), .Q(\buf [129]));
    defparam buf_129__198.GSR = "DISABLED";
    FD1S3AX buf_128__199 (.D(\buf [92]), .CK(clock), .Q(\buf [128]));
    defparam buf_128__199.GSR = "DISABLED";
    FD1S3AX buf_127__200 (.D(\buf [91]), .CK(clock), .Q(\buf [127]));
    defparam buf_127__200.GSR = "DISABLED";
    FD1S3AX buf_126__201 (.D(\buf [90]), .CK(clock), .Q(\buf [126]));
    defparam buf_126__201.GSR = "DISABLED";
    FD1S3AX buf_125__202 (.D(\buf [89]), .CK(clock), .Q(\buf [125]));
    defparam buf_125__202.GSR = "DISABLED";
    FD1S3AX buf_124__203 (.D(\buf [88]), .CK(clock), .Q(\buf [124]));
    defparam buf_124__203.GSR = "DISABLED";
    FD1S3AX buf_123__204 (.D(\buf [87]), .CK(clock), .Q(\buf [123]));
    defparam buf_123__204.GSR = "DISABLED";
    FD1S3AX buf_122__205 (.D(\buf [86]), .CK(clock), .Q(\buf [122]));
    defparam buf_122__205.GSR = "DISABLED";
    FD1S3AX buf_121__206 (.D(\buf [85]), .CK(clock), .Q(\buf [121]));
    defparam buf_121__206.GSR = "DISABLED";
    FD1S3AX buf_120__207 (.D(\buf [84]), .CK(clock), .Q(\buf [120]));
    defparam buf_120__207.GSR = "DISABLED";
    FD1S3AX buf_119__208 (.D(\buf [83]), .CK(clock), .Q(\buf [119]));
    defparam buf_119__208.GSR = "DISABLED";
    FD1S3AX buf_118__209 (.D(\buf [82]), .CK(clock), .Q(\buf [118]));
    defparam buf_118__209.GSR = "DISABLED";
    FD1S3AX buf_117__210 (.D(\buf [81]), .CK(clock), .Q(\buf [117]));
    defparam buf_117__210.GSR = "DISABLED";
    FD1S3AX buf_116__211 (.D(\buf [80]), .CK(clock), .Q(\buf [116]));
    defparam buf_116__211.GSR = "DISABLED";
    FD1S3AX buf_115__212 (.D(\buf [79]), .CK(clock), .Q(\buf [115]));
    defparam buf_115__212.GSR = "DISABLED";
    FD1S3AX buf_114__213 (.D(\buf [78]), .CK(clock), .Q(\buf [114]));
    defparam buf_114__213.GSR = "DISABLED";
    FD1S3AX buf_113__214 (.D(\buf [77]), .CK(clock), .Q(\buf [113]));
    defparam buf_113__214.GSR = "DISABLED";
    FD1S3AX buf_112__215 (.D(\buf [76]), .CK(clock), .Q(\buf [112]));
    defparam buf_112__215.GSR = "DISABLED";
    FD1S3AX buf_111__216 (.D(\buf [75]), .CK(clock), .Q(\buf [111]));
    defparam buf_111__216.GSR = "DISABLED";
    FD1S3AX buf_110__217 (.D(\buf [74]), .CK(clock), .Q(\buf [110]));
    defparam buf_110__217.GSR = "DISABLED";
    FD1S3AX buf_109__218 (.D(\buf [73]), .CK(clock), .Q(\buf [109]));
    defparam buf_109__218.GSR = "DISABLED";
    FD1S3AX buf_108__219 (.D(\buf [72]), .CK(clock), .Q(\buf [108]));
    defparam buf_108__219.GSR = "DISABLED";
    FD1S3AX buf_99__228 (.D(\buf_x[437] ), .CK(clock), .Q(\buf [99]));
    defparam buf_99__228.GSR = "DISABLED";
    FD1S3AX buf_98__229 (.D(\buf_x[436] ), .CK(clock), .Q(\buf [98]));
    defparam buf_98__229.GSR = "DISABLED";
    FD1S3AX buf_97__230 (.D(\buf_x[435] ), .CK(clock), .Q(\buf [97]));
    defparam buf_97__230.GSR = "DISABLED";
    FD1S3AX buf_96__231 (.D(\buf_x[434] ), .CK(clock), .Q(\buf [96]));
    defparam buf_96__231.GSR = "DISABLED";
    FD1S3AX buf_95__232 (.D(\buf [59]), .CK(clock), .Q(\buf [95]));
    defparam buf_95__232.GSR = "DISABLED";
    FD1S3AX buf_94__233 (.D(\buf [58]), .CK(clock), .Q(\buf [94]));
    defparam buf_94__233.GSR = "DISABLED";
    FD1S3AX buf_93__234 (.D(\buf [57]), .CK(clock), .Q(\buf [93]));
    defparam buf_93__234.GSR = "DISABLED";
    FD1S3AX buf_92__235 (.D(\buf [56]), .CK(clock), .Q(\buf [92]));
    defparam buf_92__235.GSR = "DISABLED";
    FD1S3AX buf_91__236 (.D(\buf [55]), .CK(clock), .Q(\buf [91]));
    defparam buf_91__236.GSR = "DISABLED";
    FD1S3AX buf_90__237 (.D(\buf [54]), .CK(clock), .Q(\buf [90]));
    defparam buf_90__237.GSR = "DISABLED";
    FD1S3AX buf_89__238 (.D(\buf [53]), .CK(clock), .Q(\buf [89]));
    defparam buf_89__238.GSR = "DISABLED";
    FD1S3AX buf_88__239 (.D(\buf [52]), .CK(clock), .Q(\buf [88]));
    defparam buf_88__239.GSR = "DISABLED";
    FD1S3AX buf_87__240 (.D(\buf [51]), .CK(clock), .Q(\buf [87]));
    defparam buf_87__240.GSR = "DISABLED";
    FD1S3AX buf_86__241 (.D(\buf [50]), .CK(clock), .Q(\buf [86]));
    defparam buf_86__241.GSR = "DISABLED";
    FD1S3AX buf_85__242 (.D(\buf [49]), .CK(clock), .Q(\buf [85]));
    defparam buf_85__242.GSR = "DISABLED";
    FD1S3AX buf_84__243 (.D(\buf [48]), .CK(clock), .Q(\buf [84]));
    defparam buf_84__243.GSR = "DISABLED";
    FD1S3AX buf_83__244 (.D(\buf [47]), .CK(clock), .Q(\buf [83]));
    defparam buf_83__244.GSR = "DISABLED";
    FD1S3AX buf_82__245 (.D(\buf [46]), .CK(clock), .Q(\buf [82]));
    defparam buf_82__245.GSR = "DISABLED";
    FD1S3AX buf_81__246 (.D(\buf [45]), .CK(clock), .Q(\buf [81]));
    defparam buf_81__246.GSR = "DISABLED";
    FD1S3AX buf_80__247 (.D(\buf [44]), .CK(clock), .Q(\buf [80]));
    defparam buf_80__247.GSR = "DISABLED";
    FD1S3AX buf_79__248 (.D(\buf [43]), .CK(clock), .Q(\buf [79]));
    defparam buf_79__248.GSR = "DISABLED";
    FD1S3AX buf_78__249 (.D(\buf [42]), .CK(clock), .Q(\buf [78]));
    defparam buf_78__249.GSR = "DISABLED";
    FD1S3AX buf_77__250 (.D(\buf [41]), .CK(clock), .Q(\buf [77]));
    defparam buf_77__250.GSR = "DISABLED";
    FD1S3AX buf_76__251 (.D(\buf [40]), .CK(clock), .Q(\buf [76]));
    defparam buf_76__251.GSR = "DISABLED";
    FD1S3AX buf_75__252 (.D(\buf [39]), .CK(clock), .Q(\buf [75]));
    defparam buf_75__252.GSR = "DISABLED";
    FD1S3AX buf_74__253 (.D(\buf [38]), .CK(clock), .Q(\buf [74]));
    defparam buf_74__253.GSR = "DISABLED";
    FD1S3AX buf_73__254 (.D(\buf [37]), .CK(clock), .Q(\buf [73]));
    defparam buf_73__254.GSR = "DISABLED";
    FD1S3AX buf_72__255 (.D(\buf [36]), .CK(clock), .Q(\buf [72]));
    defparam buf_72__255.GSR = "DISABLED";
    FD1S3AX buf_59__268 (.D(\nX_a1[23] ), .CK(clock), .Q(\buf [59]));
    defparam buf_59__268.GSR = "DISABLED";
    FD1S3AX buf_58__269 (.D(\nX_a1[22] ), .CK(clock), .Q(\buf [58]));
    defparam buf_58__269.GSR = "DISABLED";
    FD1S3AX buf_57__270 (.D(\nX_a1[21] ), .CK(clock), .Q(\buf [57]));
    defparam buf_57__270.GSR = "DISABLED";
    FD1S3AX buf_56__271 (.D(\nX_a1[20] ), .CK(clock), .Q(\buf [56]));
    defparam buf_56__271.GSR = "DISABLED";
    FD1S3AX buf_55__272 (.D(\nX_a1[19] ), .CK(clock), .Q(\buf [55]));
    defparam buf_55__272.GSR = "DISABLED";
    FD1S3AX buf_54__273 (.D(\nX_a1[18] ), .CK(clock), .Q(\buf [54]));
    defparam buf_54__273.GSR = "DISABLED";
    FD1S3AX buf_53__274 (.D(\nX_a1[17] ), .CK(clock), .Q(\buf [53]));
    defparam buf_53__274.GSR = "DISABLED";
    FD1S3AX buf_52__275 (.D(\nX_a1[16] ), .CK(clock), .Q(\buf [52]));
    defparam buf_52__275.GSR = "DISABLED";
    FD1S3AX buf_51__276 (.D(\nX_a1[15] ), .CK(clock), .Q(\buf [51]));
    defparam buf_51__276.GSR = "DISABLED";
    FD1S3AX buf_50__277 (.D(\nX_a1[14] ), .CK(clock), .Q(\buf [50]));
    defparam buf_50__277.GSR = "DISABLED";
    FD1S3AX buf_49__278 (.D(\nX_a1[13] ), .CK(clock), .Q(\buf [49]));
    defparam buf_49__278.GSR = "DISABLED";
    FD1S3AX buf_48__279 (.D(\nX_a1[12] ), .CK(clock), .Q(\buf [48]));
    defparam buf_48__279.GSR = "DISABLED";
    FD1S3AX buf_47__280 (.D(\nX_a1[11] ), .CK(clock), .Q(\buf [47]));
    defparam buf_47__280.GSR = "DISABLED";
    FD1S3AX buf_46__281 (.D(\nX_a1[10] ), .CK(clock), .Q(\buf [46]));
    defparam buf_46__281.GSR = "DISABLED";
    FD1S3AX buf_45__282 (.D(\nX_a1[9] ), .CK(clock), .Q(\buf [45]));
    defparam buf_45__282.GSR = "DISABLED";
    FD1S3AX buf_44__283 (.D(\nX_a1[8] ), .CK(clock), .Q(\buf [44]));
    defparam buf_44__283.GSR = "DISABLED";
    FD1S3AX buf_43__284 (.D(\nX_a1[7] ), .CK(clock), .Q(\buf [43]));
    defparam buf_43__284.GSR = "DISABLED";
    FD1S3AX buf_42__285 (.D(\nX_a1[6] ), .CK(clock), .Q(\buf [42]));
    defparam buf_42__285.GSR = "DISABLED";
    FD1S3AX buf_41__286 (.D(\nX_a1[5] ), .CK(clock), .Q(\buf [41]));
    defparam buf_41__286.GSR = "DISABLED";
    FD1S3AX buf_40__287 (.D(\nX_a1[4] ), .CK(clock), .Q(\buf [40]));
    defparam buf_40__287.GSR = "DISABLED";
    FD1S3AX buf_39__288 (.D(\nX_a1[3] ), .CK(clock), .Q(\buf [39]));
    defparam buf_39__288.GSR = "DISABLED";
    FD1S3AX buf_38__289 (.D(\nX_a1[2] ), .CK(clock), .Q(\buf [38]));
    defparam buf_38__289.GSR = "DISABLED";
    FD1S3AX buf_37__290 (.D(\nX_a1[1] ), .CK(clock), .Q(\buf [37]));
    defparam buf_37__290.GSR = "DISABLED";
    FD1S3AX buf_36__291 (.D(\nX_a1[0] ), .CK(clock), .Q(\buf [36]));
    defparam buf_36__291.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \delay(9,10) 
//

module \delay(9,10)  (\buf_r[936] , clock, \buf_x[699] , \nK_e3[7] , 
            \nK_e3[6] , \nK_e3[5] , \nK_e3[4] , \nK_e3[3] , \nK_e3[2] , 
            \nK_e3[1] , \nK_e3[0] , \buf_x[727] , \buf_x[737] , \buf_x[689] , 
            \buf_x[651] , \buf_x[661] , \buf_x[613] , \buf_x[623] );
    output \buf_r[936] ;
    input clock;
    input \buf_x[699] ;
    output \nK_e3[7] ;
    output \nK_e3[6] ;
    output \nK_e3[5] ;
    output \nK_e3[4] ;
    output \nK_e3[3] ;
    output \nK_e3[2] ;
    output \nK_e3[1] ;
    output \nK_e3[0] ;
    input \buf_x[727] ;
    input \buf_x[737] ;
    input \buf_x[689] ;
    input \buf_x[651] ;
    input \buf_x[661] ;
    input \buf_x[613] ;
    input \buf_x[623] ;
    
    wire [98:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    
    FD1S3AX buf_r_936__223 (.D(\buf_x[699] ), .CK(clock), .Q(\buf_r[936] ));
    defparam buf_r_936__223.GSR = "DISABLED";
    FD1S3AX buf_97__95 (.D(\buf [88]), .CK(clock), .Q(\nK_e3[7] ));
    defparam buf_97__95.GSR = "DISABLED";
    FD1S3AX buf_96__96 (.D(\buf [87]), .CK(clock), .Q(\nK_e3[6] ));
    defparam buf_96__96.GSR = "DISABLED";
    FD1S3AX buf_95__97 (.D(\buf [86]), .CK(clock), .Q(\nK_e3[5] ));
    defparam buf_95__97.GSR = "DISABLED";
    FD1S3AX buf_94__98 (.D(\buf [85]), .CK(clock), .Q(\nK_e3[4] ));
    defparam buf_94__98.GSR = "DISABLED";
    FD1S3AX buf_93__99 (.D(\buf [84]), .CK(clock), .Q(\nK_e3[3] ));
    defparam buf_93__99.GSR = "DISABLED";
    FD1S3AX buf_92__100 (.D(\buf [83]), .CK(clock), .Q(\nK_e3[2] ));
    defparam buf_92__100.GSR = "DISABLED";
    FD1S3AX buf_91__101 (.D(\buf [82]), .CK(clock), .Q(\nK_e3[1] ));
    defparam buf_91__101.GSR = "DISABLED";
    FD1S3AX buf_90__102 (.D(\buf [81]), .CK(clock), .Q(\nK_e3[0] ));
    defparam buf_90__102.GSR = "DISABLED";
    FD1S3AX buf_88__104 (.D(\buf [79]), .CK(clock), .Q(\buf [88]));
    defparam buf_88__104.GSR = "DISABLED";
    FD1S3AX buf_87__105 (.D(\buf [78]), .CK(clock), .Q(\buf [87]));
    defparam buf_87__105.GSR = "DISABLED";
    FD1S3AX buf_86__106 (.D(\buf [77]), .CK(clock), .Q(\buf [86]));
    defparam buf_86__106.GSR = "DISABLED";
    FD1S3AX buf_85__107 (.D(\buf [76]), .CK(clock), .Q(\buf [85]));
    defparam buf_85__107.GSR = "DISABLED";
    FD1S3AX buf_84__108 (.D(\buf [75]), .CK(clock), .Q(\buf [84]));
    defparam buf_84__108.GSR = "DISABLED";
    FD1S3AX buf_83__109 (.D(\buf [74]), .CK(clock), .Q(\buf [83]));
    defparam buf_83__109.GSR = "DISABLED";
    FD1S3AX buf_82__110 (.D(\buf [73]), .CK(clock), .Q(\buf [82]));
    defparam buf_82__110.GSR = "DISABLED";
    FD1S3AX buf_81__111 (.D(\buf [72]), .CK(clock), .Q(\buf [81]));
    defparam buf_81__111.GSR = "DISABLED";
    FD1S3AX buf_79__113 (.D(\buf [70]), .CK(clock), .Q(\buf [79]));
    defparam buf_79__113.GSR = "DISABLED";
    FD1S3AX buf_78__114 (.D(\buf [69]), .CK(clock), .Q(\buf [78]));
    defparam buf_78__114.GSR = "DISABLED";
    FD1S3AX buf_77__115 (.D(\buf [68]), .CK(clock), .Q(\buf [77]));
    defparam buf_77__115.GSR = "DISABLED";
    FD1S3AX buf_76__116 (.D(\buf [67]), .CK(clock), .Q(\buf [76]));
    defparam buf_76__116.GSR = "DISABLED";
    FD1S3AX buf_75__117 (.D(\buf [66]), .CK(clock), .Q(\buf [75]));
    defparam buf_75__117.GSR = "DISABLED";
    FD1S3AX buf_74__118 (.D(\buf [65]), .CK(clock), .Q(\buf [74]));
    defparam buf_74__118.GSR = "DISABLED";
    FD1S3AX buf_73__119 (.D(\buf [64]), .CK(clock), .Q(\buf [73]));
    defparam buf_73__119.GSR = "DISABLED";
    FD1S3AX buf_72__120 (.D(\buf [63]), .CK(clock), .Q(\buf [72]));
    defparam buf_72__120.GSR = "DISABLED";
    FD1S3AX buf_70__122 (.D(\buf [61]), .CK(clock), .Q(\buf [70]));
    defparam buf_70__122.GSR = "DISABLED";
    FD1S3AX buf_69__123 (.D(\buf [60]), .CK(clock), .Q(\buf [69]));
    defparam buf_69__123.GSR = "DISABLED";
    FD1S3AX buf_68__124 (.D(\buf [59]), .CK(clock), .Q(\buf [68]));
    defparam buf_68__124.GSR = "DISABLED";
    FD1S3AX buf_67__125 (.D(\buf [58]), .CK(clock), .Q(\buf [67]));
    defparam buf_67__125.GSR = "DISABLED";
    FD1S3AX buf_66__126 (.D(\buf [57]), .CK(clock), .Q(\buf [66]));
    defparam buf_66__126.GSR = "DISABLED";
    FD1S3AX buf_65__127 (.D(\buf [56]), .CK(clock), .Q(\buf [65]));
    defparam buf_65__127.GSR = "DISABLED";
    FD1S3AX buf_64__128 (.D(\buf [55]), .CK(clock), .Q(\buf [64]));
    defparam buf_64__128.GSR = "DISABLED";
    FD1S3AX buf_63__129 (.D(\buf [54]), .CK(clock), .Q(\buf [63]));
    defparam buf_63__129.GSR = "DISABLED";
    FD1S3AX buf_61__131 (.D(\buf [52]), .CK(clock), .Q(\buf [61]));
    defparam buf_61__131.GSR = "DISABLED";
    FD1S3AX buf_60__132 (.D(\buf [51]), .CK(clock), .Q(\buf [60]));
    defparam buf_60__132.GSR = "DISABLED";
    FD1S3AX buf_59__133 (.D(\buf [50]), .CK(clock), .Q(\buf [59]));
    defparam buf_59__133.GSR = "DISABLED";
    FD1S3AX buf_58__134 (.D(\buf [49]), .CK(clock), .Q(\buf [58]));
    defparam buf_58__134.GSR = "DISABLED";
    FD1S3AX buf_57__135 (.D(\buf [48]), .CK(clock), .Q(\buf [57]));
    defparam buf_57__135.GSR = "DISABLED";
    FD1S3AX buf_56__136 (.D(\buf [47]), .CK(clock), .Q(\buf [56]));
    defparam buf_56__136.GSR = "DISABLED";
    FD1S3AX buf_55__137 (.D(\buf [46]), .CK(clock), .Q(\buf [55]));
    defparam buf_55__137.GSR = "DISABLED";
    FD1S3AX buf_54__138 (.D(\buf [45]), .CK(clock), .Q(\buf [54]));
    defparam buf_54__138.GSR = "DISABLED";
    FD1S3AX buf_52__140 (.D(\buf [43]), .CK(clock), .Q(\buf [52]));
    defparam buf_52__140.GSR = "DISABLED";
    FD1S3AX buf_51__141 (.D(\buf [42]), .CK(clock), .Q(\buf [51]));
    defparam buf_51__141.GSR = "DISABLED";
    FD1S3AX buf_50__142 (.D(\buf [41]), .CK(clock), .Q(\buf [50]));
    defparam buf_50__142.GSR = "DISABLED";
    FD1S3AX buf_49__143 (.D(\buf [40]), .CK(clock), .Q(\buf [49]));
    defparam buf_49__143.GSR = "DISABLED";
    FD1S3AX buf_48__144 (.D(\buf [39]), .CK(clock), .Q(\buf [48]));
    defparam buf_48__144.GSR = "DISABLED";
    FD1S3AX buf_47__145 (.D(\buf [38]), .CK(clock), .Q(\buf [47]));
    defparam buf_47__145.GSR = "DISABLED";
    FD1S3AX buf_46__146 (.D(\buf [37]), .CK(clock), .Q(\buf [46]));
    defparam buf_46__146.GSR = "DISABLED";
    FD1S3AX buf_45__147 (.D(\buf [36]), .CK(clock), .Q(\buf [45]));
    defparam buf_45__147.GSR = "DISABLED";
    FD1S3AX buf_43__149 (.D(\buf [34]), .CK(clock), .Q(\buf [43]));
    defparam buf_43__149.GSR = "DISABLED";
    FD1S3AX buf_42__150 (.D(\buf [33]), .CK(clock), .Q(\buf [42]));
    defparam buf_42__150.GSR = "DISABLED";
    FD1S3AX buf_41__151 (.D(\buf [32]), .CK(clock), .Q(\buf [41]));
    defparam buf_41__151.GSR = "DISABLED";
    FD1S3AX buf_40__152 (.D(\buf [31]), .CK(clock), .Q(\buf [40]));
    defparam buf_40__152.GSR = "DISABLED";
    FD1S3AX buf_39__153 (.D(\buf [30]), .CK(clock), .Q(\buf [39]));
    defparam buf_39__153.GSR = "DISABLED";
    FD1S3AX buf_38__154 (.D(\buf [29]), .CK(clock), .Q(\buf [38]));
    defparam buf_38__154.GSR = "DISABLED";
    FD1S3AX buf_37__155 (.D(\buf [28]), .CK(clock), .Q(\buf [37]));
    defparam buf_37__155.GSR = "DISABLED";
    FD1S3AX buf_36__156 (.D(\buf [27]), .CK(clock), .Q(\buf [36]));
    defparam buf_36__156.GSR = "DISABLED";
    FD1S3AX buf_34__158 (.D(\buf [25]), .CK(clock), .Q(\buf [34]));
    defparam buf_34__158.GSR = "DISABLED";
    FD1S3AX buf_33__159 (.D(\buf [24]), .CK(clock), .Q(\buf [33]));
    defparam buf_33__159.GSR = "DISABLED";
    FD1S3AX buf_32__160 (.D(\buf [23]), .CK(clock), .Q(\buf [32]));
    defparam buf_32__160.GSR = "DISABLED";
    FD1S3AX buf_31__161 (.D(\buf [22]), .CK(clock), .Q(\buf [31]));
    defparam buf_31__161.GSR = "DISABLED";
    FD1S3AX buf_30__162 (.D(\buf [21]), .CK(clock), .Q(\buf [30]));
    defparam buf_30__162.GSR = "DISABLED";
    FD1S3AX buf_29__163 (.D(\buf [20]), .CK(clock), .Q(\buf [29]));
    defparam buf_29__163.GSR = "DISABLED";
    FD1S3AX buf_28__164 (.D(\buf [19]), .CK(clock), .Q(\buf [28]));
    defparam buf_28__164.GSR = "DISABLED";
    FD1S3AX buf_27__165 (.D(\buf [18]), .CK(clock), .Q(\buf [27]));
    defparam buf_27__165.GSR = "DISABLED";
    FD1S3AX buf_25__167 (.D(\buf [16]), .CK(clock), .Q(\buf [25]));
    defparam buf_25__167.GSR = "DISABLED";
    FD1S3AX buf_24__168 (.D(\buf [15]), .CK(clock), .Q(\buf [24]));
    defparam buf_24__168.GSR = "DISABLED";
    FD1S3AX buf_23__169 (.D(\buf [14]), .CK(clock), .Q(\buf [23]));
    defparam buf_23__169.GSR = "DISABLED";
    FD1S3AX buf_22__170 (.D(\buf_r[936] ), .CK(clock), .Q(\buf [22]));
    defparam buf_22__170.GSR = "DISABLED";
    FD1S3AX buf_21__171 (.D(\buf [12]), .CK(clock), .Q(\buf [21]));
    defparam buf_21__171.GSR = "DISABLED";
    FD1S3AX buf_20__172 (.D(\buf [11]), .CK(clock), .Q(\buf [20]));
    defparam buf_20__172.GSR = "DISABLED";
    FD1S3AX buf_19__173 (.D(\buf [10]), .CK(clock), .Q(\buf [19]));
    defparam buf_19__173.GSR = "DISABLED";
    FD1S3AX buf_18__174 (.D(\buf [9]), .CK(clock), .Q(\buf [18]));
    defparam buf_18__174.GSR = "DISABLED";
    FD1S3AX buf_16__176 (.D(\buf_x[727] ), .CK(clock), .Q(\buf [16]));
    defparam buf_16__176.GSR = "DISABLED";
    FD1S3AX buf_15__177 (.D(\buf_x[737] ), .CK(clock), .Q(\buf [15]));
    defparam buf_15__177.GSR = "DISABLED";
    FD1S3AX buf_14__178 (.D(\buf_x[689] ), .CK(clock), .Q(\buf [14]));
    defparam buf_14__178.GSR = "DISABLED";
    FD1S3AX buf_12__180 (.D(\buf_x[651] ), .CK(clock), .Q(\buf [12]));
    defparam buf_12__180.GSR = "DISABLED";
    FD1S3AX buf_11__181 (.D(\buf_x[661] ), .CK(clock), .Q(\buf [11]));
    defparam buf_11__181.GSR = "DISABLED";
    FD1S3AX buf_10__182 (.D(\buf_x[613] ), .CK(clock), .Q(\buf [10]));
    defparam buf_10__182.GSR = "DISABLED";
    FD1S3AX buf_9__183 (.D(\buf_x[623] ), .CK(clock), .Q(\buf [9]));
    defparam buf_9__183.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \delay(28,3) 
//

module \delay(28,3)  (nEY1_e1, clock, nEY1_d2);
    output [27:0]nEY1_e1;
    input clock;
    input [27:0]nEY1_d2;
    
    wire [111:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    
    FD1S3AX buf_110__89 (.D(\buf [82]), .CK(clock), .Q(nEY1_e1[26]));
    defparam buf_110__89.GSR = "DISABLED";
    FD1S3AX buf_109__90 (.D(\buf [81]), .CK(clock), .Q(nEY1_e1[25]));
    defparam buf_109__90.GSR = "DISABLED";
    FD1S3AX buf_108__91 (.D(\buf [80]), .CK(clock), .Q(nEY1_e1[24]));
    defparam buf_108__91.GSR = "DISABLED";
    FD1S3AX buf_107__92 (.D(\buf [79]), .CK(clock), .Q(nEY1_e1[23]));
    defparam buf_107__92.GSR = "DISABLED";
    FD1S3AX buf_106__93 (.D(\buf [78]), .CK(clock), .Q(nEY1_e1[22]));
    defparam buf_106__93.GSR = "DISABLED";
    FD1S3AX buf_105__94 (.D(\buf [77]), .CK(clock), .Q(nEY1_e1[21]));
    defparam buf_105__94.GSR = "DISABLED";
    FD1S3AX buf_104__95 (.D(\buf [76]), .CK(clock), .Q(nEY1_e1[20]));
    defparam buf_104__95.GSR = "DISABLED";
    FD1S3AX buf_103__96 (.D(\buf [75]), .CK(clock), .Q(nEY1_e1[19]));
    defparam buf_103__96.GSR = "DISABLED";
    FD1S3AX buf_102__97 (.D(\buf [74]), .CK(clock), .Q(nEY1_e1[18]));
    defparam buf_102__97.GSR = "DISABLED";
    FD1S3AX buf_101__98 (.D(\buf [73]), .CK(clock), .Q(nEY1_e1[17]));
    defparam buf_101__98.GSR = "DISABLED";
    FD1S3AX buf_100__99 (.D(\buf [72]), .CK(clock), .Q(nEY1_e1[16]));
    defparam buf_100__99.GSR = "DISABLED";
    FD1S3AX buf_99__100 (.D(\buf [71]), .CK(clock), .Q(nEY1_e1[15]));
    defparam buf_99__100.GSR = "DISABLED";
    FD1S3AX buf_98__101 (.D(\buf [70]), .CK(clock), .Q(nEY1_e1[14]));
    defparam buf_98__101.GSR = "DISABLED";
    FD1S3AX buf_97__102 (.D(\buf [69]), .CK(clock), .Q(nEY1_e1[13]));
    defparam buf_97__102.GSR = "DISABLED";
    FD1S3AX buf_96__103 (.D(\buf [68]), .CK(clock), .Q(nEY1_e1[12]));
    defparam buf_96__103.GSR = "DISABLED";
    FD1S3AX buf_95__104 (.D(\buf [67]), .CK(clock), .Q(nEY1_e1[11]));
    defparam buf_95__104.GSR = "DISABLED";
    FD1S3AX buf_94__105 (.D(\buf [66]), .CK(clock), .Q(nEY1_e1[10]));
    defparam buf_94__105.GSR = "DISABLED";
    FD1S3AX buf_93__106 (.D(\buf [65]), .CK(clock), .Q(nEY1_e1[9]));
    defparam buf_93__106.GSR = "DISABLED";
    FD1S3AX buf_92__107 (.D(\buf [64]), .CK(clock), .Q(nEY1_e1[8]));
    defparam buf_92__107.GSR = "DISABLED";
    FD1S3AX buf_91__108 (.D(\buf [63]), .CK(clock), .Q(nEY1_e1[7]));
    defparam buf_91__108.GSR = "DISABLED";
    FD1S3AX buf_90__109 (.D(\buf [62]), .CK(clock), .Q(nEY1_e1[6]));
    defparam buf_90__109.GSR = "DISABLED";
    FD1S3AX buf_89__110 (.D(\buf [61]), .CK(clock), .Q(nEY1_e1[5]));
    defparam buf_89__110.GSR = "DISABLED";
    FD1S3AX buf_88__111 (.D(\buf [60]), .CK(clock), .Q(nEY1_e1[4]));
    defparam buf_88__111.GSR = "DISABLED";
    FD1S3AX buf_87__112 (.D(\buf [59]), .CK(clock), .Q(nEY1_e1[3]));
    defparam buf_87__112.GSR = "DISABLED";
    FD1S3AX buf_86__113 (.D(\buf [58]), .CK(clock), .Q(nEY1_e1[2]));
    defparam buf_86__113.GSR = "DISABLED";
    FD1S3AX buf_85__114 (.D(\buf [57]), .CK(clock), .Q(nEY1_e1[1]));
    defparam buf_85__114.GSR = "DISABLED";
    FD1S3AX buf_84__115 (.D(\buf [56]), .CK(clock), .Q(nEY1_e1[0]));
    defparam buf_84__115.GSR = "DISABLED";
    FD1S3AX buf_83__116 (.D(\buf [55]), .CK(clock), .Q(\buf [83]));
    defparam buf_83__116.GSR = "DISABLED";
    FD1S3AX buf_82__117 (.D(\buf [54]), .CK(clock), .Q(\buf [82]));
    defparam buf_82__117.GSR = "DISABLED";
    FD1S3AX buf_81__118 (.D(\buf [53]), .CK(clock), .Q(\buf [81]));
    defparam buf_81__118.GSR = "DISABLED";
    FD1S3AX buf_80__119 (.D(\buf [52]), .CK(clock), .Q(\buf [80]));
    defparam buf_80__119.GSR = "DISABLED";
    FD1S3AX buf_79__120 (.D(\buf [51]), .CK(clock), .Q(\buf [79]));
    defparam buf_79__120.GSR = "DISABLED";
    FD1S3AX buf_78__121 (.D(\buf [50]), .CK(clock), .Q(\buf [78]));
    defparam buf_78__121.GSR = "DISABLED";
    FD1S3AX buf_77__122 (.D(\buf [49]), .CK(clock), .Q(\buf [77]));
    defparam buf_77__122.GSR = "DISABLED";
    FD1S3AX buf_76__123 (.D(\buf [48]), .CK(clock), .Q(\buf [76]));
    defparam buf_76__123.GSR = "DISABLED";
    FD1S3AX buf_75__124 (.D(\buf [47]), .CK(clock), .Q(\buf [75]));
    defparam buf_75__124.GSR = "DISABLED";
    FD1S3AX buf_74__125 (.D(\buf [46]), .CK(clock), .Q(\buf [74]));
    defparam buf_74__125.GSR = "DISABLED";
    FD1S3AX buf_73__126 (.D(\buf [45]), .CK(clock), .Q(\buf [73]));
    defparam buf_73__126.GSR = "DISABLED";
    FD1S3AX buf_72__127 (.D(\buf [44]), .CK(clock), .Q(\buf [72]));
    defparam buf_72__127.GSR = "DISABLED";
    FD1S3AX buf_71__128 (.D(\buf [43]), .CK(clock), .Q(\buf [71]));
    defparam buf_71__128.GSR = "DISABLED";
    FD1S3AX buf_70__129 (.D(\buf [42]), .CK(clock), .Q(\buf [70]));
    defparam buf_70__129.GSR = "DISABLED";
    FD1S3AX buf_69__130 (.D(\buf [41]), .CK(clock), .Q(\buf [69]));
    defparam buf_69__130.GSR = "DISABLED";
    FD1S3AX buf_68__131 (.D(\buf [40]), .CK(clock), .Q(\buf [68]));
    defparam buf_68__131.GSR = "DISABLED";
    FD1S3AX buf_67__132 (.D(\buf [39]), .CK(clock), .Q(\buf [67]));
    defparam buf_67__132.GSR = "DISABLED";
    FD1S3AX buf_66__133 (.D(\buf [38]), .CK(clock), .Q(\buf [66]));
    defparam buf_66__133.GSR = "DISABLED";
    FD1S3AX buf_65__134 (.D(\buf [37]), .CK(clock), .Q(\buf [65]));
    defparam buf_65__134.GSR = "DISABLED";
    FD1S3AX buf_64__135 (.D(\buf [36]), .CK(clock), .Q(\buf [64]));
    defparam buf_64__135.GSR = "DISABLED";
    FD1S3AX buf_63__136 (.D(\buf [35]), .CK(clock), .Q(\buf [63]));
    defparam buf_63__136.GSR = "DISABLED";
    FD1S3AX buf_62__137 (.D(\buf [34]), .CK(clock), .Q(\buf [62]));
    defparam buf_62__137.GSR = "DISABLED";
    FD1S3AX buf_61__138 (.D(\buf [33]), .CK(clock), .Q(\buf [61]));
    defparam buf_61__138.GSR = "DISABLED";
    FD1S3AX buf_60__139 (.D(\buf [32]), .CK(clock), .Q(\buf [60]));
    defparam buf_60__139.GSR = "DISABLED";
    FD1S3AX buf_59__140 (.D(\buf [31]), .CK(clock), .Q(\buf [59]));
    defparam buf_59__140.GSR = "DISABLED";
    FD1S3AX buf_58__141 (.D(\buf [30]), .CK(clock), .Q(\buf [58]));
    defparam buf_58__141.GSR = "DISABLED";
    FD1S3AX buf_57__142 (.D(\buf [29]), .CK(clock), .Q(\buf [57]));
    defparam buf_57__142.GSR = "DISABLED";
    FD1S3AX buf_56__143 (.D(\buf [28]), .CK(clock), .Q(\buf [56]));
    defparam buf_56__143.GSR = "DISABLED";
    FD1S3AX buf_55__144 (.D(nEY1_d2[27]), .CK(clock), .Q(\buf [55]));
    defparam buf_55__144.GSR = "DISABLED";
    FD1S3AX buf_54__145 (.D(nEY1_d2[26]), .CK(clock), .Q(\buf [54]));
    defparam buf_54__145.GSR = "DISABLED";
    FD1S3AX buf_53__146 (.D(nEY1_d2[25]), .CK(clock), .Q(\buf [53]));
    defparam buf_53__146.GSR = "DISABLED";
    FD1S3AX buf_52__147 (.D(nEY1_d2[24]), .CK(clock), .Q(\buf [52]));
    defparam buf_52__147.GSR = "DISABLED";
    FD1S3AX buf_51__148 (.D(nEY1_d2[23]), .CK(clock), .Q(\buf [51]));
    defparam buf_51__148.GSR = "DISABLED";
    FD1S3AX buf_50__149 (.D(nEY1_d2[22]), .CK(clock), .Q(\buf [50]));
    defparam buf_50__149.GSR = "DISABLED";
    FD1S3AX buf_49__150 (.D(nEY1_d2[21]), .CK(clock), .Q(\buf [49]));
    defparam buf_49__150.GSR = "DISABLED";
    FD1S3AX buf_48__151 (.D(nEY1_d2[20]), .CK(clock), .Q(\buf [48]));
    defparam buf_48__151.GSR = "DISABLED";
    FD1S3AX buf_47__152 (.D(nEY1_d2[19]), .CK(clock), .Q(\buf [47]));
    defparam buf_47__152.GSR = "DISABLED";
    FD1S3AX buf_46__153 (.D(nEY1_d2[18]), .CK(clock), .Q(\buf [46]));
    defparam buf_46__153.GSR = "DISABLED";
    FD1S3AX buf_45__154 (.D(nEY1_d2[17]), .CK(clock), .Q(\buf [45]));
    defparam buf_45__154.GSR = "DISABLED";
    FD1S3AX buf_44__155 (.D(nEY1_d2[16]), .CK(clock), .Q(\buf [44]));
    defparam buf_44__155.GSR = "DISABLED";
    FD1S3AX buf_43__156 (.D(nEY1_d2[15]), .CK(clock), .Q(\buf [43]));
    defparam buf_43__156.GSR = "DISABLED";
    FD1S3AX buf_42__157 (.D(nEY1_d2[14]), .CK(clock), .Q(\buf [42]));
    defparam buf_42__157.GSR = "DISABLED";
    FD1S3AX buf_41__158 (.D(nEY1_d2[13]), .CK(clock), .Q(\buf [41]));
    defparam buf_41__158.GSR = "DISABLED";
    FD1S3AX buf_40__159 (.D(nEY1_d2[12]), .CK(clock), .Q(\buf [40]));
    defparam buf_40__159.GSR = "DISABLED";
    FD1S3AX buf_39__160 (.D(nEY1_d2[11]), .CK(clock), .Q(\buf [39]));
    defparam buf_39__160.GSR = "DISABLED";
    FD1S3AX buf_38__161 (.D(nEY1_d2[10]), .CK(clock), .Q(\buf [38]));
    defparam buf_38__161.GSR = "DISABLED";
    FD1S3AX buf_37__162 (.D(nEY1_d2[9]), .CK(clock), .Q(\buf [37]));
    defparam buf_37__162.GSR = "DISABLED";
    FD1S3AX buf_36__163 (.D(nEY1_d2[8]), .CK(clock), .Q(\buf [36]));
    defparam buf_36__163.GSR = "DISABLED";
    FD1S3AX buf_35__164 (.D(nEY1_d2[7]), .CK(clock), .Q(\buf [35]));
    defparam buf_35__164.GSR = "DISABLED";
    FD1S3AX buf_34__165 (.D(nEY1_d2[6]), .CK(clock), .Q(\buf [34]));
    defparam buf_34__165.GSR = "DISABLED";
    FD1S3AX buf_33__166 (.D(nEY1_d2[5]), .CK(clock), .Q(\buf [33]));
    defparam buf_33__166.GSR = "DISABLED";
    FD1S3AX buf_32__167 (.D(nEY1_d2[4]), .CK(clock), .Q(\buf [32]));
    defparam buf_32__167.GSR = "DISABLED";
    FD1S3AX buf_31__168 (.D(nEY1_d2[3]), .CK(clock), .Q(\buf [31]));
    defparam buf_31__168.GSR = "DISABLED";
    FD1S3AX buf_30__169 (.D(nEY1_d2[2]), .CK(clock), .Q(\buf [30]));
    defparam buf_30__169.GSR = "DISABLED";
    FD1S3AX buf_29__170 (.D(nEY1_d2[1]), .CK(clock), .Q(\buf [29]));
    defparam buf_29__170.GSR = "DISABLED";
    FD1S3AX buf_28__171 (.D(nEY1_d2[0]), .CK(clock), .Q(\buf [28]));
    defparam buf_28__171.GSR = "DISABLED";
    FD1S3AX buf_111__88 (.D(\buf [83]), .CK(clock), .Q(nEY1_e1[27]));
    defparam buf_111__88.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \delay(28,3)_U25 
//

module \delay(28,3)_U25  (nEY1_d2, clock, \nEY1_c1[24] , \nEY1_c1[23] , 
            \nEY1_c1[22] , \nEY1_c1[21] , \nEY1_c1[20] , \nEY1_c1[19] , 
            \nEY1_c1[18] , \nEY1_c1[17] , \nEY1_c1[16] , \nEY1_c1[15] , 
            \nEY1_c1[14] , \nEY1_c1[13] , \nEY1_c1[12] , \nEY1_c1[11] , 
            \nEY1_c1[10] , \nEY1_c1[9] , \nEY1_c1[8] , \nEY1_c1[7] , 
            \nEY1_c1[6] , \nEY1_c1[5] , \nEY1_c1[4] , \nEY1_c1[3] , 
            \nEY1_c1[2] , \nEY1_c1[1] , \nEY1_c1[0] , \nY1_c1[7] , \nY_c1[27] , 
            n62787, \nEY1_c1[25] );
    output [27:0]nEY1_d2;
    input clock;
    input \nEY1_c1[24] ;
    input \nEY1_c1[23] ;
    input \nEY1_c1[22] ;
    input \nEY1_c1[21] ;
    input \nEY1_c1[20] ;
    input \nEY1_c1[19] ;
    input \nEY1_c1[18] ;
    input \nEY1_c1[17] ;
    input \nEY1_c1[16] ;
    input \nEY1_c1[15] ;
    input \nEY1_c1[14] ;
    input \nEY1_c1[13] ;
    input \nEY1_c1[12] ;
    input \nEY1_c1[11] ;
    input \nEY1_c1[10] ;
    input \nEY1_c1[9] ;
    input \nEY1_c1[8] ;
    input \nEY1_c1[7] ;
    input \nEY1_c1[6] ;
    input \nEY1_c1[5] ;
    input \nEY1_c1[4] ;
    input \nEY1_c1[3] ;
    input \nEY1_c1[2] ;
    input \nEY1_c1[1] ;
    input \nEY1_c1[0] ;
    input \nY1_c1[7] ;
    input \nY_c1[27] ;
    input n62787;
    input \nEY1_c1[25] ;
    
    wire [111:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    
    FD1S3AX buf_110__89 (.D(\buf [82]), .CK(clock), .Q(nEY1_d2[26]));
    defparam buf_110__89.GSR = "DISABLED";
    FD1S3AX buf_109__90 (.D(\buf [81]), .CK(clock), .Q(nEY1_d2[25]));
    defparam buf_109__90.GSR = "DISABLED";
    FD1S3AX buf_108__91 (.D(\buf [80]), .CK(clock), .Q(nEY1_d2[24]));
    defparam buf_108__91.GSR = "DISABLED";
    FD1S3AX buf_107__92 (.D(\buf [79]), .CK(clock), .Q(nEY1_d2[23]));
    defparam buf_107__92.GSR = "DISABLED";
    FD1S3AX buf_106__93 (.D(\buf [78]), .CK(clock), .Q(nEY1_d2[22]));
    defparam buf_106__93.GSR = "DISABLED";
    FD1S3AX buf_105__94 (.D(\buf [77]), .CK(clock), .Q(nEY1_d2[21]));
    defparam buf_105__94.GSR = "DISABLED";
    FD1S3AX buf_104__95 (.D(\buf [76]), .CK(clock), .Q(nEY1_d2[20]));
    defparam buf_104__95.GSR = "DISABLED";
    FD1S3AX buf_103__96 (.D(\buf [75]), .CK(clock), .Q(nEY1_d2[19]));
    defparam buf_103__96.GSR = "DISABLED";
    FD1S3AX buf_102__97 (.D(\buf [74]), .CK(clock), .Q(nEY1_d2[18]));
    defparam buf_102__97.GSR = "DISABLED";
    FD1S3AX buf_101__98 (.D(\buf [73]), .CK(clock), .Q(nEY1_d2[17]));
    defparam buf_101__98.GSR = "DISABLED";
    FD1S3AX buf_100__99 (.D(\buf [72]), .CK(clock), .Q(nEY1_d2[16]));
    defparam buf_100__99.GSR = "DISABLED";
    FD1S3AX buf_99__100 (.D(\buf [71]), .CK(clock), .Q(nEY1_d2[15]));
    defparam buf_99__100.GSR = "DISABLED";
    FD1S3AX buf_98__101 (.D(\buf [70]), .CK(clock), .Q(nEY1_d2[14]));
    defparam buf_98__101.GSR = "DISABLED";
    FD1S3AX buf_97__102 (.D(\buf [69]), .CK(clock), .Q(nEY1_d2[13]));
    defparam buf_97__102.GSR = "DISABLED";
    FD1S3AX buf_96__103 (.D(\buf [68]), .CK(clock), .Q(nEY1_d2[12]));
    defparam buf_96__103.GSR = "DISABLED";
    FD1S3AX buf_95__104 (.D(\buf [67]), .CK(clock), .Q(nEY1_d2[11]));
    defparam buf_95__104.GSR = "DISABLED";
    FD1S3AX buf_94__105 (.D(\buf [66]), .CK(clock), .Q(nEY1_d2[10]));
    defparam buf_94__105.GSR = "DISABLED";
    FD1S3AX buf_93__106 (.D(\buf [65]), .CK(clock), .Q(nEY1_d2[9]));
    defparam buf_93__106.GSR = "DISABLED";
    FD1S3AX buf_92__107 (.D(\buf [64]), .CK(clock), .Q(nEY1_d2[8]));
    defparam buf_92__107.GSR = "DISABLED";
    FD1S3AX buf_91__108 (.D(\buf [63]), .CK(clock), .Q(nEY1_d2[7]));
    defparam buf_91__108.GSR = "DISABLED";
    FD1S3AX buf_90__109 (.D(\buf [62]), .CK(clock), .Q(nEY1_d2[6]));
    defparam buf_90__109.GSR = "DISABLED";
    FD1S3AX buf_89__110 (.D(\buf [61]), .CK(clock), .Q(nEY1_d2[5]));
    defparam buf_89__110.GSR = "DISABLED";
    FD1S3AX buf_88__111 (.D(\buf [60]), .CK(clock), .Q(nEY1_d2[4]));
    defparam buf_88__111.GSR = "DISABLED";
    FD1S3AX buf_87__112 (.D(\buf [59]), .CK(clock), .Q(nEY1_d2[3]));
    defparam buf_87__112.GSR = "DISABLED";
    FD1S3AX buf_86__113 (.D(\buf [58]), .CK(clock), .Q(nEY1_d2[2]));
    defparam buf_86__113.GSR = "DISABLED";
    FD1S3AX buf_85__114 (.D(\buf [57]), .CK(clock), .Q(nEY1_d2[1]));
    defparam buf_85__114.GSR = "DISABLED";
    FD1S3AX buf_84__115 (.D(\buf [56]), .CK(clock), .Q(nEY1_d2[0]));
    defparam buf_84__115.GSR = "DISABLED";
    FD1S3AX buf_83__116 (.D(\buf [55]), .CK(clock), .Q(\buf [83]));
    defparam buf_83__116.GSR = "DISABLED";
    FD1S3AX buf_82__117 (.D(\buf [54]), .CK(clock), .Q(\buf [82]));
    defparam buf_82__117.GSR = "DISABLED";
    FD1S3AX buf_81__118 (.D(\buf [53]), .CK(clock), .Q(\buf [81]));
    defparam buf_81__118.GSR = "DISABLED";
    FD1S3AX buf_80__119 (.D(\nEY1_c1[24] ), .CK(clock), .Q(\buf [80]));
    defparam buf_80__119.GSR = "DISABLED";
    FD1S3AX buf_79__120 (.D(\nEY1_c1[23] ), .CK(clock), .Q(\buf [79]));
    defparam buf_79__120.GSR = "DISABLED";
    FD1S3AX buf_78__121 (.D(\nEY1_c1[22] ), .CK(clock), .Q(\buf [78]));
    defparam buf_78__121.GSR = "DISABLED";
    FD1S3AX buf_77__122 (.D(\nEY1_c1[21] ), .CK(clock), .Q(\buf [77]));
    defparam buf_77__122.GSR = "DISABLED";
    FD1S3AX buf_76__123 (.D(\nEY1_c1[20] ), .CK(clock), .Q(\buf [76]));
    defparam buf_76__123.GSR = "DISABLED";
    FD1S3AX buf_75__124 (.D(\nEY1_c1[19] ), .CK(clock), .Q(\buf [75]));
    defparam buf_75__124.GSR = "DISABLED";
    FD1S3AX buf_74__125 (.D(\nEY1_c1[18] ), .CK(clock), .Q(\buf [74]));
    defparam buf_74__125.GSR = "DISABLED";
    FD1S3AX buf_73__126 (.D(\nEY1_c1[17] ), .CK(clock), .Q(\buf [73]));
    defparam buf_73__126.GSR = "DISABLED";
    FD1S3AX buf_72__127 (.D(\nEY1_c1[16] ), .CK(clock), .Q(\buf [72]));
    defparam buf_72__127.GSR = "DISABLED";
    FD1S3AX buf_71__128 (.D(\nEY1_c1[15] ), .CK(clock), .Q(\buf [71]));
    defparam buf_71__128.GSR = "DISABLED";
    FD1S3AX buf_70__129 (.D(\nEY1_c1[14] ), .CK(clock), .Q(\buf [70]));
    defparam buf_70__129.GSR = "DISABLED";
    FD1S3AX buf_69__130 (.D(\nEY1_c1[13] ), .CK(clock), .Q(\buf [69]));
    defparam buf_69__130.GSR = "DISABLED";
    FD1S3AX buf_68__131 (.D(\nEY1_c1[12] ), .CK(clock), .Q(\buf [68]));
    defparam buf_68__131.GSR = "DISABLED";
    FD1S3AX buf_67__132 (.D(\nEY1_c1[11] ), .CK(clock), .Q(\buf [67]));
    defparam buf_67__132.GSR = "DISABLED";
    FD1S3AX buf_66__133 (.D(\nEY1_c1[10] ), .CK(clock), .Q(\buf [66]));
    defparam buf_66__133.GSR = "DISABLED";
    FD1S3AX buf_65__134 (.D(\nEY1_c1[9] ), .CK(clock), .Q(\buf [65]));
    defparam buf_65__134.GSR = "DISABLED";
    FD1S3AX buf_64__135 (.D(\nEY1_c1[8] ), .CK(clock), .Q(\buf [64]));
    defparam buf_64__135.GSR = "DISABLED";
    FD1S3AX buf_63__136 (.D(\nEY1_c1[7] ), .CK(clock), .Q(\buf [63]));
    defparam buf_63__136.GSR = "DISABLED";
    FD1S3AX buf_62__137 (.D(\nEY1_c1[6] ), .CK(clock), .Q(\buf [62]));
    defparam buf_62__137.GSR = "DISABLED";
    FD1S3AX buf_61__138 (.D(\nEY1_c1[5] ), .CK(clock), .Q(\buf [61]));
    defparam buf_61__138.GSR = "DISABLED";
    FD1S3AX buf_60__139 (.D(\nEY1_c1[4] ), .CK(clock), .Q(\buf [60]));
    defparam buf_60__139.GSR = "DISABLED";
    FD1S3AX buf_59__140 (.D(\nEY1_c1[3] ), .CK(clock), .Q(\buf [59]));
    defparam buf_59__140.GSR = "DISABLED";
    FD1S3AX buf_58__141 (.D(\nEY1_c1[2] ), .CK(clock), .Q(\buf [58]));
    defparam buf_58__141.GSR = "DISABLED";
    FD1S3AX buf_57__142 (.D(\nEY1_c1[1] ), .CK(clock), .Q(\buf [57]));
    defparam buf_57__142.GSR = "DISABLED";
    FD1S3AX buf_56__143 (.D(\nEY1_c1[0] ), .CK(clock), .Q(\buf [56]));
    defparam buf_56__143.GSR = "DISABLED";
    FD1S3AX buf_55__144 (.D(\nY1_c1[7] ), .CK(clock), .Q(\buf [55]));
    defparam buf_55__144.GSR = "DISABLED";
    FD1S3JX buf_54__145 (.D(n62787), .CK(clock), .PD(\nY_c1[27] ), .Q(\buf [54]));
    defparam buf_54__145.GSR = "DISABLED";
    FD1S3AX buf_53__146 (.D(\nEY1_c1[25] ), .CK(clock), .Q(\buf [53]));
    defparam buf_53__146.GSR = "DISABLED";
    FD1S3AX buf_111__88 (.D(\buf [83]), .CK(clock), .Q(nEY1_d2[27]));
    defparam buf_111__88.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \delay(34,14) 
//

module \delay(34,14)  (\buf[474] , clock, \exp_a[32] );
    output \buf[474] ;
    input clock;
    input \exp_a[32] ;
    
    wire [509:0]\buf ;   // c:/users/yisong/documents/new/mlp/fp_exp.vhd(286[10:13])
    
    FD1S3AX buf_474__515 (.D(\buf [440]), .CK(clock), .Q(\buf[474] ));
    defparam buf_474__515.GSR = "DISABLED";
    FD1S3AX buf_440__549 (.D(\buf [406]), .CK(clock), .Q(\buf [440]));
    defparam buf_440__549.GSR = "DISABLED";
    FD1S3AX buf_406__583 (.D(\buf [372]), .CK(clock), .Q(\buf [406]));
    defparam buf_406__583.GSR = "DISABLED";
    FD1S3AX buf_372__617 (.D(\buf [338]), .CK(clock), .Q(\buf [372]));
    defparam buf_372__617.GSR = "DISABLED";
    FD1S3AX buf_338__651 (.D(\buf [304]), .CK(clock), .Q(\buf [338]));
    defparam buf_338__651.GSR = "DISABLED";
    FD1S3AX buf_304__685 (.D(\buf [270]), .CK(clock), .Q(\buf [304]));
    defparam buf_304__685.GSR = "DISABLED";
    FD1S3AX buf_270__719 (.D(\buf [236]), .CK(clock), .Q(\buf [270]));
    defparam buf_270__719.GSR = "DISABLED";
    FD1S3AX buf_236__753 (.D(\buf [202]), .CK(clock), .Q(\buf [236]));
    defparam buf_236__753.GSR = "DISABLED";
    FD1S3AX buf_202__787 (.D(\buf [168]), .CK(clock), .Q(\buf [202]));
    defparam buf_202__787.GSR = "DISABLED";
    FD1S3AX buf_168__821 (.D(\buf [134]), .CK(clock), .Q(\buf [168]));
    defparam buf_168__821.GSR = "DISABLED";
    FD1S3AX buf_134__855 (.D(\buf [100]), .CK(clock), .Q(\buf [134]));
    defparam buf_134__855.GSR = "DISABLED";
    FD1S3AX buf_100__889 (.D(\buf [66]), .CK(clock), .Q(\buf [100]));
    defparam buf_100__889.GSR = "DISABLED";
    FD1S3AX buf_66__923 (.D(\exp_a[32] ), .CK(clock), .Q(\buf [66]));
    defparam buf_66__923.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \fp_div(32,24,8) 
//

module \fp_div(32,24,8)  (GND_net, clock, n73815, alu_b, alu_a, div_c, 
            div_ce, n73814);
    input GND_net;
    input clock;
    input n73815;
    input [31:0]alu_b;
    input [31:0]alu_a;
    output [31:0]div_c;
    input div_ce;
    input n73814;
    
    wire [31:0]B_int;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(59[18:23])
    wire [31:0]A_int;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(59[11:16])
    wire [8:0]exp_Biased;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(66[23:33])
    wire [26:0]\QQ_in[1] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[25] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[26] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[24] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[22] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[23] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[20] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[21] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[18] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[19] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[16] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[17] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[14] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[15] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[12] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[13] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[10] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[11] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [8:0]exp_Biased_Norm;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(66[35:50])
    wire [26:0]\QQ_in[6] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[7] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[8] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [31:0]FP_Z_int;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(59[25:33])
    wire [26:0]\QQ_in[9] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[4] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[5] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[2] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire [26:0]\QQ_in[3] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(44[11:16])
    wire expB_FF;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(64[20:27])
    wire expA_FF;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(64[11:18])
    
    wire n61603, n17202, n416, n17200;
    wire [22:0]n10674;
    
    wire n61604, n61602, n17206, n17204, n61601, n17210, n17208, 
        n61600, n17214, n17212, n61599, n17218, n17216, n61598, 
        n17222, n17220, n61597, n17226, n17224, n61596, n17230, 
        n17228, n61595, n17234, n17232, n17, n15, n61593;
    wire [8:0]n14;
    wire [8:0]n284;
    
    wire n61592, n61591, n61590, n417, n70750, n10, n70745, n423, 
        n70754, n424, n70753, n418, n70752, n422, n70751, n421, 
        n420, n70749, n419, n70748, n28, n38, n24, n36, n42, 
        n32, n40, n44, n31, n66210, n28_adj_447, n38_adj_448, 
        n24_adj_449, n36_adj_450, n42_adj_451, n32_adj_452, n40_adj_453, 
        n44_adj_454, n31_adj_455, n22395, n10_adj_456, n1, n24032, 
        n21749, n10_adj_457, n66951, n66953, n16_adj_458, n11, n21, 
        n15_adj_459;
    wire [31:0]n65;
    
    wire n61536, n61535, n61534, n61533, n66694, n415, n17196, 
        n17198, n17192, n17194, n10_adj_460, n14_adj_461, n10_adj_462, 
        n14_adj_463, n16_adj_464, n15_adj_465, n4, n9256, n61605;
    
    CCU2D add_3814_19 (.A0(n17202), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17200), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61603), 
          .COUT(n61604), .S0(n10674[17]), .S1(n10674[18]));
    defparam add_3814_19.INIT0 = 16'he111;
    defparam add_3814_19.INIT1 = 16'he111;
    defparam add_3814_19.INJECT1_0 = "NO";
    defparam add_3814_19.INJECT1_1 = "NO";
    FD1P3AX B_int_i0_i0 (.D(alu_b[0]), .SP(n73815), .CK(clock), .Q(B_int[0]));
    defparam B_int_i0_i0.GSR = "DISABLED";
    FD1P3AX A_int_i0_i0 (.D(alu_a[0]), .SP(n73815), .CK(clock), .Q(A_int[0]));
    defparam A_int_i0_i0.GSR = "DISABLED";
    CCU2D add_3814_17 (.A0(n17206), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17204), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61602), 
          .COUT(n61603), .S0(n10674[15]), .S1(n10674[16]));
    defparam add_3814_17.INIT0 = 16'he111;
    defparam add_3814_17.INIT1 = 16'he111;
    defparam add_3814_17.INJECT1_0 = "NO";
    defparam add_3814_17.INJECT1_1 = "NO";
    CCU2D add_3814_15 (.A0(n17210), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17208), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61601), 
          .COUT(n61602), .S0(n10674[13]), .S1(n10674[14]));
    defparam add_3814_15.INIT0 = 16'he111;
    defparam add_3814_15.INIT1 = 16'he111;
    defparam add_3814_15.INJECT1_0 = "NO";
    defparam add_3814_15.INJECT1_1 = "NO";
    CCU2D add_3814_13 (.A0(n17214), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17212), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61600), 
          .COUT(n61601), .S0(n10674[11]), .S1(n10674[12]));
    defparam add_3814_13.INIT0 = 16'he111;
    defparam add_3814_13.INIT1 = 16'he111;
    defparam add_3814_13.INJECT1_0 = "NO";
    defparam add_3814_13.INJECT1_1 = "NO";
    CCU2D add_3814_11 (.A0(n17218), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17216), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61599), 
          .COUT(n61600), .S0(n10674[9]), .S1(n10674[10]));
    defparam add_3814_11.INIT0 = 16'he111;
    defparam add_3814_11.INIT1 = 16'he111;
    defparam add_3814_11.INJECT1_0 = "NO";
    defparam add_3814_11.INJECT1_1 = "NO";
    CCU2D add_3814_9 (.A0(n17222), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17220), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61598), 
          .COUT(n61599), .S0(n10674[7]), .S1(n10674[8]));
    defparam add_3814_9.INIT0 = 16'he111;
    defparam add_3814_9.INIT1 = 16'he111;
    defparam add_3814_9.INJECT1_0 = "NO";
    defparam add_3814_9.INJECT1_1 = "NO";
    CCU2D add_3814_7 (.A0(n17226), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17224), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61597), 
          .COUT(n61598), .S0(n10674[5]), .S1(n10674[6]));
    defparam add_3814_7.INIT0 = 16'he111;
    defparam add_3814_7.INIT1 = 16'he111;
    defparam add_3814_7.INJECT1_0 = "NO";
    defparam add_3814_7.INJECT1_1 = "NO";
    CCU2D add_3814_5 (.A0(n17230), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17228), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61596), 
          .COUT(n61597), .S0(n10674[3]), .S1(n10674[4]));
    defparam add_3814_5.INIT0 = 16'he111;
    defparam add_3814_5.INIT1 = 16'he111;
    defparam add_3814_5.INJECT1_0 = "NO";
    defparam add_3814_5.INJECT1_1 = "NO";
    CCU2D add_3814_3 (.A0(n17234), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17232), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61595), 
          .COUT(n61596), .S0(n10674[1]), .S1(n10674[2]));
    defparam add_3814_3.INIT0 = 16'he111;
    defparam add_3814_3.INIT1 = 16'he111;
    defparam add_3814_3.INJECT1_0 = "NO";
    defparam add_3814_3.INJECT1_1 = "NO";
    CCU2D add_3814_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n416), .B1(n17), .C1(n15), .D1(GND_net), .COUT(n61595), 
          .S1(n10674[0]));
    defparam add_3814_1.INIT0 = 16'hF000;
    defparam add_3814_1.INIT1 = 16'he414;
    defparam add_3814_1.INJECT1_0 = "NO";
    defparam add_3814_1.INJECT1_1 = "NO";
    CCU2D add_31_9 (.A0(n14[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n14[8]), .B1(n14[7]), .C1(GND_net), .D1(GND_net), .CIN(n61593), 
          .S0(n284[7]), .S1(n284[8]));
    defparam add_31_9.INIT0 = 16'haaaa;
    defparam add_31_9.INIT1 = 16'h9999;
    defparam add_31_9.INJECT1_0 = "NO";
    defparam add_31_9.INJECT1_1 = "NO";
    CCU2D add_31_7 (.A0(exp_Biased[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_Biased[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61592), .COUT(n61593), .S0(n284[5]), .S1(n284[6]));
    defparam add_31_7.INIT0 = 16'h5555;
    defparam add_31_7.INIT1 = 16'h5555;
    defparam add_31_7.INJECT1_0 = "NO";
    defparam add_31_7.INJECT1_1 = "NO";
    CCU2D add_31_5 (.A0(exp_Biased[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_Biased[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61591), .COUT(n61592), .S0(n284[3]), .S1(n284[4]));
    defparam add_31_5.INIT0 = 16'h5555;
    defparam add_31_5.INIT1 = 16'h5555;
    defparam add_31_5.INJECT1_0 = "NO";
    defparam add_31_5.INJECT1_1 = "NO";
    CCU2D add_31_3 (.A0(exp_Biased[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_Biased[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61590), .COUT(n61591), .S0(n284[1]), .S1(n284[2]));
    defparam add_31_3.INIT0 = 16'h5555;
    defparam add_31_3.INIT1 = 16'h5555;
    defparam add_31_3.INJECT1_0 = "NO";
    defparam add_31_3.INJECT1_1 = "NO";
    LUT4 i27786_2_lut_4_lut_4_lut (.A(n14[7]), .B(n416), .C(\QQ_in[1] [0]), 
         .D(n284[7]), .Z(n417)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!((D)+!C)))) */ ;
    defparam i27786_2_lut_4_lut_4_lut.init = 16'h3101;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n14[7]), .B(n70750), .C(\QQ_in[1] [0]), 
         .D(n284[7]), .Z(n10)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'hc404;
    LUT4 mux_33_i8_3_lut_rep_775_3_lut (.A(n14[7]), .B(\QQ_in[1] [0]), .C(n284[7]), 
         .Z(n70745)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_33_i8_3_lut_rep_775_3_lut.init = 16'hd1d1;
    CCU2D add_31_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(exp_Biased[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n61590), .S1(n284[0]));
    defparam add_31_1.INIT0 = 16'hF000;
    defparam add_31_1.INIT1 = 16'h5555;
    defparam add_31_1.INJECT1_0 = "NO";
    defparam add_31_1.INJECT1_1 = "NO";
    LUT4 i13602_3_lut (.A(\QQ_in[25] [24]), .B(\QQ_in[26] [25]), .C(\QQ_in[1] [0]), 
         .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13602_3_lut.init = 16'hcaca;
    LUT4 i13606_3_lut (.A(\QQ_in[24] [23]), .B(\QQ_in[25] [24]), .C(\QQ_in[1] [0]), 
         .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13606_3_lut.init = 16'hcaca;
    LUT4 mux_156_i6_3_lut (.A(\QQ_in[22] [21]), .B(\QQ_in[23] [22]), .C(\QQ_in[1] [0]), 
         .Z(n17232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i6_3_lut.init = 16'hcaca;
    LUT4 mux_156_i5_3_lut (.A(\QQ_in[23] [22]), .B(\QQ_in[24] [23]), .C(\QQ_in[1] [0]), 
         .Z(n17234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i5_3_lut.init = 16'hcaca;
    LUT4 mux_156_i8_3_lut (.A(\QQ_in[20] [19]), .B(\QQ_in[21] [20]), .C(\QQ_in[1] [0]), 
         .Z(n17228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i8_3_lut.init = 16'hcaca;
    LUT4 mux_156_i7_3_lut (.A(\QQ_in[21] [20]), .B(\QQ_in[22] [21]), .C(\QQ_in[1] [0]), 
         .Z(n17230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i7_3_lut.init = 16'hcaca;
    LUT4 mux_156_i10_3_lut (.A(\QQ_in[18] [17]), .B(\QQ_in[19] [18]), .C(\QQ_in[1] [0]), 
         .Z(n17224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i10_3_lut.init = 16'hcaca;
    LUT4 mux_156_i9_3_lut (.A(\QQ_in[19] [18]), .B(\QQ_in[20] [19]), .C(\QQ_in[1] [0]), 
         .Z(n17226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i9_3_lut.init = 16'hcaca;
    LUT4 mux_156_i12_3_lut (.A(\QQ_in[16] [15]), .B(\QQ_in[17] [16]), .C(\QQ_in[1] [0]), 
         .Z(n17220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i12_3_lut.init = 16'hcaca;
    LUT4 mux_156_i11_3_lut (.A(\QQ_in[17] [16]), .B(\QQ_in[18] [17]), .C(\QQ_in[1] [0]), 
         .Z(n17222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i11_3_lut.init = 16'hcaca;
    LUT4 mux_156_i14_3_lut (.A(\QQ_in[14] [13]), .B(\QQ_in[15] [14]), .C(\QQ_in[1] [0]), 
         .Z(n17216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i14_3_lut.init = 16'hcaca;
    LUT4 mux_156_i13_3_lut (.A(\QQ_in[15] [14]), .B(\QQ_in[16] [15]), .C(\QQ_in[1] [0]), 
         .Z(n17218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i13_3_lut.init = 16'hcaca;
    LUT4 mux_156_i16_3_lut (.A(\QQ_in[12] [11]), .B(\QQ_in[13] [12]), .C(\QQ_in[1] [0]), 
         .Z(n17212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i16_3_lut.init = 16'hcaca;
    LUT4 mux_156_i15_3_lut (.A(\QQ_in[13] [12]), .B(\QQ_in[14] [13]), .C(\QQ_in[1] [0]), 
         .Z(n17214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i15_3_lut.init = 16'hcaca;
    LUT4 mux_156_i18_3_lut (.A(\QQ_in[10] [9]), .B(\QQ_in[11] [10]), .C(\QQ_in[1] [0]), 
         .Z(n17208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i18_3_lut.init = 16'hcaca;
    LUT4 mux_156_i17_3_lut (.A(\QQ_in[11] [10]), .B(\QQ_in[12] [11]), .C(\QQ_in[1] [0]), 
         .Z(n17210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i17_3_lut.init = 16'hcaca;
    LUT4 i27792_2_lut_4_lut (.A(exp_Biased[1]), .B(n284[1]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n423)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27792_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i2_3_lut_rep_784 (.A(exp_Biased[1]), .B(n284[1]), .C(\QQ_in[1] [0]), 
         .Z(n70754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i2_3_lut_rep_784.init = 16'hcaca;
    LUT4 i27793_2_lut_4_lut (.A(exp_Biased[0]), .B(n284[0]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n424)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27793_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i1_3_lut_rep_783 (.A(exp_Biased[0]), .B(n284[0]), .C(\QQ_in[1] [0]), 
         .Z(n70753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i1_3_lut_rep_783.init = 16'hcaca;
    LUT4 i27787_2_lut_4_lut (.A(exp_Biased[6]), .B(n284[6]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n418)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27787_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i7_3_lut_rep_782 (.A(exp_Biased[6]), .B(n284[6]), .C(\QQ_in[1] [0]), 
         .Z(n70752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i7_3_lut_rep_782.init = 16'hcaca;
    LUT4 i27791_2_lut_4_lut (.A(exp_Biased[2]), .B(n284[2]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n422)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27791_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i3_3_lut_rep_781 (.A(exp_Biased[2]), .B(n284[2]), .C(\QQ_in[1] [0]), 
         .Z(n70751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i3_3_lut_rep_781.init = 16'hcaca;
    LUT4 i27790_2_lut_4_lut (.A(exp_Biased[3]), .B(n284[3]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n421)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27790_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i4_3_lut_rep_780 (.A(exp_Biased[3]), .B(n284[3]), .C(\QQ_in[1] [0]), 
         .Z(n70750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i4_3_lut_rep_780.init = 16'hcaca;
    LUT4 i27789_2_lut_4_lut (.A(exp_Biased[4]), .B(n284[4]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n420)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27789_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i5_3_lut_rep_779 (.A(exp_Biased[4]), .B(n284[4]), .C(\QQ_in[1] [0]), 
         .Z(n70749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i5_3_lut_rep_779.init = 16'hcaca;
    LUT4 i27788_2_lut_4_lut (.A(exp_Biased[5]), .B(n284[5]), .C(\QQ_in[1] [0]), 
         .D(n416), .Z(n419)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i27788_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_33_i6_3_lut_rep_778 (.A(exp_Biased[5]), .B(n284[5]), .C(\QQ_in[1] [0]), 
         .Z(n70748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_33_i6_3_lut_rep_778.init = 16'hcaca;
    LUT4 mux_33_i9_4_lut (.A(n14[8]), .B(n284[8]), .C(\QQ_in[1] [0]), 
         .D(n14[7]), .Z(exp_Biased_Norm[8])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_33_i9_4_lut.init = 16'hc5ca;
    LUT4 i5_2_lut (.A(A_int[12]), .B(A_int[10]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i15_4_lut (.A(A_int[18]), .B(A_int[3]), .C(A_int[11]), .D(A_int[22]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(A_int[19]), .B(A_int[0]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i13_4_lut (.A(A_int[17]), .B(A_int[6]), .C(A_int[5]), .D(A_int[16]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(A_int[4]), .B(n38), .C(n28), .D(A_int[14]), .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(A_int[15]), .B(A_int[21]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(A_int[7]), .B(A_int[2]), .C(A_int[1]), .D(A_int[20]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(A_int[9]), .B(n42), .C(n36), .D(n24), .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(A_int[13]), .B(A_int[8]), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(n31), .B(n44), .C(n40), .D(n32), .Z(n66210)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut_adj_815 (.A(B_int[6]), .B(B_int[10]), .Z(n28_adj_447)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut_adj_815.init = 16'heeee;
    LUT4 i15_4_lut_adj_816 (.A(B_int[13]), .B(B_int[16]), .C(B_int[9]), 
         .D(B_int[17]), .Z(n38_adj_448)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_816.init = 16'hfffe;
    LUT4 i1_2_lut_adj_817 (.A(B_int[21]), .B(B_int[14]), .Z(n24_adj_449)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_817.init = 16'heeee;
    LUT4 i13_4_lut_adj_818 (.A(B_int[12]), .B(B_int[20]), .C(B_int[18]), 
         .D(B_int[19]), .Z(n36_adj_450)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_818.init = 16'hfffe;
    LUT4 i19_4_lut_adj_819 (.A(B_int[15]), .B(n38_adj_448), .C(n28_adj_447), 
         .D(B_int[5]), .Z(n42_adj_451)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_819.init = 16'hfffe;
    LUT4 i9_2_lut_adj_820 (.A(B_int[0]), .B(B_int[22]), .Z(n32_adj_452)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut_adj_820.init = 16'heeee;
    LUT4 i17_4_lut_adj_821 (.A(B_int[4]), .B(B_int[11]), .C(B_int[8]), 
         .D(B_int[1]), .Z(n40_adj_453)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_821.init = 16'hfffe;
    LUT4 i21_4_lut_adj_822 (.A(B_int[2]), .B(n42_adj_451), .C(n36_adj_450), 
         .D(n24_adj_449), .Z(n44_adj_454)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut_adj_822.init = 16'hfffe;
    LUT4 i8_2_lut_adj_823 (.A(B_int[3]), .B(B_int[7]), .Z(n31_adj_455)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut_adj_823.init = 16'heeee;
    LUT4 i22_4_lut_adj_824 (.A(n31_adj_455), .B(n44_adj_454), .C(n40_adj_453), 
         .D(n32_adj_452), .Z(n22395)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut_adj_824.init = 16'hfffe;
    LUT4 i2_2_lut (.A(B_int[25]), .B(B_int[27]), .Z(n10_adj_456)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i6_4_lut (.A(B_int[26]), .B(B_int[24]), .C(B_int[28]), .D(B_int[30]), 
         .Z(n1)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    FD1P3IX FP_Z_i0_i1 (.D(n10674[1]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[1]));
    defparam FP_Z_i0_i1.GSR = "DISABLED";
    LUT4 i7_4_lut (.A(B_int[23]), .B(n1), .C(n10_adj_456), .D(B_int[29]), 
         .Z(n21749)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 mux_156_i22_3_lut (.A(\QQ_in[6] [5]), .B(\QQ_in[7] [6]), .C(\QQ_in[1] [0]), 
         .Z(n17200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i22_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_825 (.A(A_int[25]), .B(A_int[26]), .Z(n10_adj_457)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_825.init = 16'heeee;
    LUT4 i54043_4_lut (.A(n70751), .B(n70750), .C(n70749), .D(n70748), 
         .Z(n66951)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54043_4_lut.init = 16'hfffe;
    LUT4 i54045_3_lut (.A(n70754), .B(n70753), .C(n70752), .Z(n66953)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i54045_3_lut.init = 16'hfefe;
    LUT4 i7_4_lut_adj_826 (.A(A_int[27]), .B(n66210), .C(A_int[23]), .D(n10_adj_457), 
         .Z(n16_adj_458)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_826.init = 16'hfffe;
    LUT4 i1_2_lut_adj_827 (.A(n21749), .B(n22395), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_827.init = 16'heeee;
    LUT4 i21_4_lut_adj_828 (.A(n66953), .B(exp_Biased_Norm[8]), .C(n70745), 
         .D(n66951), .Z(n21)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i21_4_lut_adj_828.init = 16'hc0c5;
    LUT4 i6_4_lut_adj_829 (.A(A_int[29]), .B(A_int[30]), .C(A_int[24]), 
         .D(A_int[28]), .Z(n15_adj_459)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_829.init = 16'hfffe;
    LUT4 i1_4_lut (.A(n15_adj_459), .B(n21), .C(n11), .D(n16_adj_458), 
         .Z(n416)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'hccdc;
    LUT4 mux_156_i21_3_lut (.A(\QQ_in[7] [6]), .B(\QQ_in[8] [7]), .C(\QQ_in[1] [0]), 
         .Z(n17202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i21_3_lut.init = 16'hcaca;
    FD1P3AX A_int_i0_i30 (.D(alu_a[30]), .SP(n73815), .CK(clock), .Q(A_int[30]));
    defparam A_int_i0_i30.GSR = "DISABLED";
    FD1P3AX A_int_i0_i29 (.D(alu_a[29]), .SP(n73815), .CK(clock), .Q(A_int[29]));
    defparam A_int_i0_i29.GSR = "DISABLED";
    FD1P3AX A_int_i0_i28 (.D(alu_a[28]), .SP(n73815), .CK(clock), .Q(A_int[28]));
    defparam A_int_i0_i28.GSR = "DISABLED";
    FD1P3AX A_int_i0_i27 (.D(alu_a[27]), .SP(n73815), .CK(clock), .Q(A_int[27]));
    defparam A_int_i0_i27.GSR = "DISABLED";
    FD1P3AX A_int_i0_i26 (.D(alu_a[26]), .SP(n73815), .CK(clock), .Q(A_int[26]));
    defparam A_int_i0_i26.GSR = "DISABLED";
    FD1P3AX A_int_i0_i25 (.D(alu_a[25]), .SP(n73815), .CK(clock), .Q(A_int[25]));
    defparam A_int_i0_i25.GSR = "DISABLED";
    FD1P3AX A_int_i0_i24 (.D(alu_a[24]), .SP(n73815), .CK(clock), .Q(A_int[24]));
    defparam A_int_i0_i24.GSR = "DISABLED";
    FD1P3AX A_int_i0_i23 (.D(alu_a[23]), .SP(n73815), .CK(clock), .Q(A_int[23]));
    defparam A_int_i0_i23.GSR = "DISABLED";
    FD1P3AX A_int_i0_i22 (.D(alu_a[22]), .SP(n73815), .CK(clock), .Q(A_int[22]));
    defparam A_int_i0_i22.GSR = "DISABLED";
    FD1P3AX A_int_i0_i21 (.D(alu_a[21]), .SP(n73815), .CK(clock), .Q(A_int[21]));
    defparam A_int_i0_i21.GSR = "DISABLED";
    FD1P3AX A_int_i0_i20 (.D(alu_a[20]), .SP(n73815), .CK(clock), .Q(A_int[20]));
    defparam A_int_i0_i20.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i2 (.D(n10674[2]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[2]));
    defparam FP_Z_i0_i2.GSR = "DISABLED";
    FD1P3AX A_int_i0_i19 (.D(alu_a[19]), .SP(n73815), .CK(clock), .Q(A_int[19]));
    defparam A_int_i0_i19.GSR = "DISABLED";
    FD1P3AX A_int_i0_i18 (.D(alu_a[18]), .SP(n73815), .CK(clock), .Q(A_int[18]));
    defparam A_int_i0_i18.GSR = "DISABLED";
    FD1P3AX A_int_i0_i17 (.D(alu_a[17]), .SP(n73815), .CK(clock), .Q(A_int[17]));
    defparam A_int_i0_i17.GSR = "DISABLED";
    FD1P3AX A_int_i0_i16 (.D(alu_a[16]), .SP(n73815), .CK(clock), .Q(A_int[16]));
    defparam A_int_i0_i16.GSR = "DISABLED";
    FD1P3AX A_int_i0_i15 (.D(alu_a[15]), .SP(n73815), .CK(clock), .Q(A_int[15]));
    defparam A_int_i0_i15.GSR = "DISABLED";
    FD1P3AX A_int_i0_i14 (.D(alu_a[14]), .SP(n73815), .CK(clock), .Q(A_int[14]));
    defparam A_int_i0_i14.GSR = "DISABLED";
    FD1P3AX A_int_i0_i13 (.D(alu_a[13]), .SP(n73815), .CK(clock), .Q(A_int[13]));
    defparam A_int_i0_i13.GSR = "DISABLED";
    FD1P3AX A_int_i0_i12 (.D(alu_a[12]), .SP(n73815), .CK(clock), .Q(A_int[12]));
    defparam A_int_i0_i12.GSR = "DISABLED";
    FD1P3AX A_int_i0_i11 (.D(alu_a[11]), .SP(n73815), .CK(clock), .Q(A_int[11]));
    defparam A_int_i0_i11.GSR = "DISABLED";
    FD1P3AX A_int_i0_i10 (.D(alu_a[10]), .SP(n73815), .CK(clock), .Q(A_int[10]));
    defparam A_int_i0_i10.GSR = "DISABLED";
    FD1P3AX A_int_i0_i9 (.D(alu_a[9]), .SP(n73815), .CK(clock), .Q(A_int[9]));
    defparam A_int_i0_i9.GSR = "DISABLED";
    FD1P3AX A_int_i0_i8 (.D(alu_a[8]), .SP(n73815), .CK(clock), .Q(A_int[8]));
    defparam A_int_i0_i8.GSR = "DISABLED";
    FD1P3AX A_int_i0_i7 (.D(alu_a[7]), .SP(n73815), .CK(clock), .Q(A_int[7]));
    defparam A_int_i0_i7.GSR = "DISABLED";
    FD1P3AX A_int_i0_i6 (.D(alu_a[6]), .SP(n73815), .CK(clock), .Q(A_int[6]));
    defparam A_int_i0_i6.GSR = "DISABLED";
    FD1P3AX A_int_i0_i5 (.D(alu_a[5]), .SP(n73815), .CK(clock), .Q(A_int[5]));
    defparam A_int_i0_i5.GSR = "DISABLED";
    FD1P3AX A_int_i0_i4 (.D(alu_a[4]), .SP(n73815), .CK(clock), .Q(A_int[4]));
    defparam A_int_i0_i4.GSR = "DISABLED";
    FD1P3AX A_int_i0_i3 (.D(alu_a[3]), .SP(n73815), .CK(clock), .Q(A_int[3]));
    defparam A_int_i0_i3.GSR = "DISABLED";
    FD1P3AX A_int_i0_i2 (.D(alu_a[2]), .SP(n73815), .CK(clock), .Q(A_int[2]));
    defparam A_int_i0_i2.GSR = "DISABLED";
    FD1P3AX A_int_i0_i1 (.D(alu_a[1]), .SP(n73815), .CK(clock), .Q(A_int[1]));
    defparam A_int_i0_i1.GSR = "DISABLED";
    FD1P3AX FP_Z_i0_i31 (.D(FP_Z_int[31]), .SP(n73815), .CK(clock), .Q(div_c[31]));
    defparam FP_Z_i0_i31.GSR = "DISABLED";
    FD1P3AX FP_Z_i0_i22 (.D(FP_Z_int[22]), .SP(n73815), .CK(clock), .Q(div_c[22]));
    defparam FP_Z_i0_i22.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i3 (.D(n10674[3]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[3]));
    defparam FP_Z_i0_i3.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i4 (.D(n10674[4]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[4]));
    defparam FP_Z_i0_i4.GSR = "DISABLED";
    FD1P3AX B_int_i0_i31 (.D(alu_b[31]), .SP(div_ce), .CK(clock), .Q(B_int[31]));
    defparam B_int_i0_i31.GSR = "DISABLED";
    FD1P3AX B_int_i0_i30 (.D(alu_b[30]), .SP(div_ce), .CK(clock), .Q(B_int[30]));
    defparam B_int_i0_i30.GSR = "DISABLED";
    FD1P3AX B_int_i0_i29 (.D(alu_b[29]), .SP(div_ce), .CK(clock), .Q(B_int[29]));
    defparam B_int_i0_i29.GSR = "DISABLED";
    FD1P3AX B_int_i0_i28 (.D(alu_b[28]), .SP(div_ce), .CK(clock), .Q(B_int[28]));
    defparam B_int_i0_i28.GSR = "DISABLED";
    FD1P3AX B_int_i0_i27 (.D(alu_b[27]), .SP(div_ce), .CK(clock), .Q(B_int[27]));
    defparam B_int_i0_i27.GSR = "DISABLED";
    FD1P3AX B_int_i0_i26 (.D(alu_b[26]), .SP(div_ce), .CK(clock), .Q(B_int[26]));
    defparam B_int_i0_i26.GSR = "DISABLED";
    FD1P3AX B_int_i0_i25 (.D(alu_b[25]), .SP(div_ce), .CK(clock), .Q(B_int[25]));
    defparam B_int_i0_i25.GSR = "DISABLED";
    FD1P3AX B_int_i0_i24 (.D(alu_b[24]), .SP(div_ce), .CK(clock), .Q(B_int[24]));
    defparam B_int_i0_i24.GSR = "DISABLED";
    FD1P3AX B_int_i0_i23 (.D(alu_b[23]), .SP(div_ce), .CK(clock), .Q(B_int[23]));
    defparam B_int_i0_i23.GSR = "DISABLED";
    FD1P3AX B_int_i0_i22 (.D(alu_b[22]), .SP(div_ce), .CK(clock), .Q(B_int[22]));
    defparam B_int_i0_i22.GSR = "DISABLED";
    FD1P3AX B_int_i0_i21 (.D(alu_b[21]), .SP(div_ce), .CK(clock), .Q(B_int[21]));
    defparam B_int_i0_i21.GSR = "DISABLED";
    FD1P3AX B_int_i0_i20 (.D(alu_b[20]), .SP(div_ce), .CK(clock), .Q(B_int[20]));
    defparam B_int_i0_i20.GSR = "DISABLED";
    FD1P3AX B_int_i0_i19 (.D(alu_b[19]), .SP(div_ce), .CK(clock), .Q(B_int[19]));
    defparam B_int_i0_i19.GSR = "DISABLED";
    FD1P3AX B_int_i0_i18 (.D(alu_b[18]), .SP(div_ce), .CK(clock), .Q(B_int[18]));
    defparam B_int_i0_i18.GSR = "DISABLED";
    FD1P3AX B_int_i0_i17 (.D(alu_b[17]), .SP(div_ce), .CK(clock), .Q(B_int[17]));
    defparam B_int_i0_i17.GSR = "DISABLED";
    FD1P3AX B_int_i0_i16 (.D(alu_b[16]), .SP(div_ce), .CK(clock), .Q(B_int[16]));
    defparam B_int_i0_i16.GSR = "DISABLED";
    FD1P3AX B_int_i0_i15 (.D(alu_b[15]), .SP(div_ce), .CK(clock), .Q(B_int[15]));
    defparam B_int_i0_i15.GSR = "DISABLED";
    FD1P3AX B_int_i0_i14 (.D(alu_b[14]), .SP(div_ce), .CK(clock), .Q(B_int[14]));
    defparam B_int_i0_i14.GSR = "DISABLED";
    FD1P3AX B_int_i0_i13 (.D(alu_b[13]), .SP(div_ce), .CK(clock), .Q(B_int[13]));
    defparam B_int_i0_i13.GSR = "DISABLED";
    FD1P3AX B_int_i0_i12 (.D(alu_b[12]), .SP(div_ce), .CK(clock), .Q(B_int[12]));
    defparam B_int_i0_i12.GSR = "DISABLED";
    FD1P3AX B_int_i0_i11 (.D(alu_b[11]), .SP(div_ce), .CK(clock), .Q(B_int[11]));
    defparam B_int_i0_i11.GSR = "DISABLED";
    FD1P3AX B_int_i0_i10 (.D(alu_b[10]), .SP(div_ce), .CK(clock), .Q(B_int[10]));
    defparam B_int_i0_i10.GSR = "DISABLED";
    FD1P3AX B_int_i0_i9 (.D(alu_b[9]), .SP(div_ce), .CK(clock), .Q(B_int[9]));
    defparam B_int_i0_i9.GSR = "DISABLED";
    FD1P3AX B_int_i0_i8 (.D(alu_b[8]), .SP(div_ce), .CK(clock), .Q(B_int[8]));
    defparam B_int_i0_i8.GSR = "DISABLED";
    FD1P3AX B_int_i0_i7 (.D(alu_b[7]), .SP(div_ce), .CK(clock), .Q(B_int[7]));
    defparam B_int_i0_i7.GSR = "DISABLED";
    FD1P3AX B_int_i0_i6 (.D(alu_b[6]), .SP(div_ce), .CK(clock), .Q(B_int[6]));
    defparam B_int_i0_i6.GSR = "DISABLED";
    FD1P3AX B_int_i0_i5 (.D(alu_b[5]), .SP(div_ce), .CK(clock), .Q(B_int[5]));
    defparam B_int_i0_i5.GSR = "DISABLED";
    FD1P3AX B_int_i0_i4 (.D(alu_b[4]), .SP(div_ce), .CK(clock), .Q(B_int[4]));
    defparam B_int_i0_i4.GSR = "DISABLED";
    FD1P3AX B_int_i0_i3 (.D(alu_b[3]), .SP(div_ce), .CK(clock), .Q(B_int[3]));
    defparam B_int_i0_i3.GSR = "DISABLED";
    FD1P3AX B_int_i0_i2 (.D(alu_b[2]), .SP(div_ce), .CK(clock), .Q(B_int[2]));
    defparam B_int_i0_i2.GSR = "DISABLED";
    FD1P3AX B_int_i0_i1 (.D(alu_b[1]), .SP(div_ce), .CK(clock), .Q(B_int[1]));
    defparam B_int_i0_i1.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i5 (.D(n10674[5]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[5]));
    defparam FP_Z_i0_i5.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i6 (.D(n10674[6]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[6]));
    defparam FP_Z_i0_i6.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i7 (.D(n10674[7]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[7]));
    defparam FP_Z_i0_i7.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i8 (.D(n10674[8]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[8]));
    defparam FP_Z_i0_i8.GSR = "DISABLED";
    LUT4 mux_156_i20_3_lut (.A(\QQ_in[8] [7]), .B(\QQ_in[9] [8]), .C(\QQ_in[1] [0]), 
         .Z(n17204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i20_3_lut.init = 16'hcaca;
    LUT4 mux_156_i19_3_lut (.A(\QQ_in[9] [8]), .B(\QQ_in[10] [9]), .C(\QQ_in[1] [0]), 
         .Z(n17206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i19_3_lut.init = 16'hcaca;
    FD1P3AX A_int_rep_3__i31 (.D(alu_a[31]), .SP(div_ce), .CK(clock), 
            .Q(n65[31]));
    defparam A_int_rep_3__i31.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i9 (.D(n10674[9]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[9]));
    defparam FP_Z_i0_i9.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i10 (.D(n10674[10]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[10]));
    defparam FP_Z_i0_i10.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i11 (.D(n10674[11]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[11]));
    defparam FP_Z_i0_i11.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i12 (.D(n10674[12]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[12]));
    defparam FP_Z_i0_i12.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i13 (.D(n10674[13]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[13]));
    defparam FP_Z_i0_i13.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i14 (.D(n10674[14]), .SP(div_ce), .CD(n24032), .CK(clock), 
            .Q(div_c[14]));
    defparam FP_Z_i0_i14.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i15 (.D(n10674[15]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[15]));
    defparam FP_Z_i0_i15.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i16 (.D(n10674[16]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[16]));
    defparam FP_Z_i0_i16.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i17 (.D(n10674[17]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[17]));
    defparam FP_Z_i0_i17.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i18 (.D(n10674[18]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[18]));
    defparam FP_Z_i0_i18.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i19 (.D(n10674[19]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[19]));
    defparam FP_Z_i0_i19.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i20 (.D(n10674[20]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[20]));
    defparam FP_Z_i0_i20.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i21 (.D(n10674[21]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[21]));
    defparam FP_Z_i0_i21.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i23 (.D(n424), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[23]));
    defparam FP_Z_i0_i23.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i24 (.D(n423), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[24]));
    defparam FP_Z_i0_i24.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i25 (.D(n422), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[25]));
    defparam FP_Z_i0_i25.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i26 (.D(n421), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[26]));
    defparam FP_Z_i0_i26.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i27 (.D(n420), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[27]));
    defparam FP_Z_i0_i27.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i28 (.D(n419), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[28]));
    defparam FP_Z_i0_i28.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i29 (.D(n418), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[29]));
    defparam FP_Z_i0_i29.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i30 (.D(n417), .SP(n73815), .PD(n24032), .CK(clock), 
            .Q(div_c[30]));
    defparam FP_Z_i0_i30.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i0 (.D(n10674[0]), .SP(n73815), .CD(n24032), .CK(clock), 
            .Q(div_c[0]));
    defparam FP_Z_i0_i0.GSR = "DISABLED";
    CCU2D add_49663_add_2_9 (.A0(B_int[30]), .B0(A_int[30]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61536), .S0(n14[7]), .S1(n14[8]));
    defparam add_49663_add_2_9.INIT0 = 16'ha999;
    defparam add_49663_add_2_9.INIT1 = 16'h0fff;
    defparam add_49663_add_2_9.INJECT1_0 = "NO";
    defparam add_49663_add_2_9.INJECT1_1 = "NO";
    CCU2D add_49663_add_2_7 (.A0(B_int[28]), .B0(A_int[28]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[29]), .B1(A_int[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61535), .COUT(n61536), .S0(exp_Biased[5]), 
          .S1(exp_Biased[6]));
    defparam add_49663_add_2_7.INIT0 = 16'ha999;
    defparam add_49663_add_2_7.INIT1 = 16'ha999;
    defparam add_49663_add_2_7.INJECT1_0 = "NO";
    defparam add_49663_add_2_7.INJECT1_1 = "NO";
    CCU2D add_49663_add_2_5 (.A0(B_int[26]), .B0(A_int[26]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[27]), .B1(A_int[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61534), .COUT(n61535), .S0(exp_Biased[3]), 
          .S1(exp_Biased[4]));
    defparam add_49663_add_2_5.INIT0 = 16'ha999;
    defparam add_49663_add_2_5.INIT1 = 16'ha999;
    defparam add_49663_add_2_5.INJECT1_0 = "NO";
    defparam add_49663_add_2_5.INJECT1_1 = "NO";
    CCU2D add_49663_add_2_3 (.A0(B_int[24]), .B0(A_int[24]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[25]), .B1(A_int[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61533), .COUT(n61534), .S0(exp_Biased[1]), 
          .S1(exp_Biased[2]));
    defparam add_49663_add_2_3.INIT0 = 16'ha999;
    defparam add_49663_add_2_3.INIT1 = 16'ha999;
    defparam add_49663_add_2_3.INJECT1_0 = "NO";
    defparam add_49663_add_2_3.INJECT1_1 = "NO";
    CCU2D add_49663_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[23]), .B1(A_int[23]), .C1(GND_net), 
          .D1(GND_net), .COUT(n61533), .S1(exp_Biased[0]));
    defparam add_49663_add_2_1.INIT0 = 16'hF000;
    defparam add_49663_add_2_1.INIT1 = 16'ha999;
    defparam add_49663_add_2_1.INJECT1_0 = "NO";
    defparam add_49663_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(n10674[22]), .B(n66694), .C(n415), .Z(FP_Z_int[22])) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i1_3_lut.init = 16'hcece;
    LUT4 i27_2_lut (.A(n65[31]), .B(B_int[31]), .Z(FP_Z_int[31])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i27_2_lut.init = 16'h6666;
    LUT4 mux_156_i24_3_lut (.A(\QQ_in[4] [3]), .B(\QQ_in[5] [4]), .C(\QQ_in[1] [0]), 
         .Z(n17196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i24_3_lut.init = 16'hcaca;
    LUT4 mux_156_i23_3_lut (.A(\QQ_in[5] [4]), .B(\QQ_in[6] [5]), .C(\QQ_in[1] [0]), 
         .Z(n17198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i23_3_lut.init = 16'hcaca;
    LUT4 mux_156_i26_3_lut (.A(\QQ_in[2] [1]), .B(\QQ_in[3] [2]), .C(\QQ_in[1] [0]), 
         .Z(n17192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i26_3_lut.init = 16'hcaca;
    LUT4 mux_156_i25_3_lut (.A(\QQ_in[3] [2]), .B(\QQ_in[4] [3]), .C(\QQ_in[1] [0]), 
         .Z(n17194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_156_i25_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_adj_830 (.A(B_int[25]), .B(B_int[27]), .Z(n10_adj_460)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_830.init = 16'h8888;
    LUT4 i6_4_lut_adj_831 (.A(B_int[26]), .B(B_int[24]), .C(B_int[28]), 
         .D(B_int[30]), .Z(n14_adj_461)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_831.init = 16'h8000;
    LUT4 i7_4_lut_adj_832 (.A(B_int[23]), .B(n14_adj_461), .C(n10_adj_460), 
         .D(B_int[29]), .Z(expB_FF)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_832.init = 16'h8000;
    LUT4 i2_2_lut_adj_833 (.A(A_int[27]), .B(A_int[24]), .Z(n10_adj_462)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_833.init = 16'h8888;
    LUT4 i6_4_lut_adj_834 (.A(A_int[26]), .B(A_int[23]), .C(A_int[28]), 
         .D(A_int[30]), .Z(n14_adj_463)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_834.init = 16'h8000;
    LUT4 i7_4_lut_adj_835 (.A(A_int[25]), .B(n14_adj_463), .C(n10_adj_462), 
         .D(A_int[29]), .Z(expA_FF)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_835.init = 16'h8000;
    LUT4 i1_4_lut_adj_836 (.A(expA_FF), .B(expB_FF), .C(n66210), .D(n22395), 
         .Z(n66694)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_836.init = 16'heca0;
    LUT4 i7_4_lut_adj_837 (.A(n70754), .B(n70748), .C(n70749), .D(n10), 
         .Z(n16_adj_464)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_837.init = 16'h8000;
    LUT4 i6_4_lut_adj_838 (.A(n70751), .B(exp_Biased_Norm[8]), .C(n70753), 
         .D(n70752), .Z(n15_adj_465)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i6_4_lut_adj_838.init = 16'h2000;
    LUT4 i1_4_lut_adj_839 (.A(n15_adj_465), .B(n70745), .C(n16_adj_464), 
         .D(exp_Biased_Norm[8]), .Z(n4)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut_adj_839.init = 16'hb3a0;
    LUT4 i2_4_lut (.A(n21749), .B(expA_FF), .C(n4), .D(expB_FF), .Z(n415)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hfffd;
    LUT4 i12369_3_lut (.A(n73814), .B(n415), .C(n66694), .Z(n24032)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i12369_3_lut.init = 16'ha8a8;
    LUT4 i3063_1_lut (.A(\QQ_in[1] [0]), .Z(n9256)) /* synthesis lut_function=(!(A)) */ ;
    defparam i3063_1_lut.init = 16'h5555;
    CCU2D add_3814_23 (.A0(n17194), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17192), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61605), 
          .S0(n10674[21]), .S1(n10674[22]));
    defparam add_3814_23.INIT0 = 16'he111;
    defparam add_3814_23.INIT1 = 16'he111;
    defparam add_3814_23.INJECT1_0 = "NO";
    defparam add_3814_23.INJECT1_1 = "NO";
    CCU2D add_3814_21 (.A0(n17198), .B0(n416), .C0(GND_net), .D0(GND_net), 
          .A1(n17196), .B1(n416), .C1(GND_net), .D1(GND_net), .CIN(n61604), 
          .COUT(n61605), .S0(n10674[19]), .S1(n10674[20]));
    defparam add_3814_21.INIT0 = 16'he111;
    defparam add_3814_21.INIT1 = 16'he111;
    defparam add_3814_21.INJECT1_0 = "NO";
    defparam add_3814_21.INJECT1_1 = "NO";
    \div_nr_wsticky(24,27)  a_div (.\QQ_in[22][21] (\QQ_in[22] [21]), .\QQ_in[21][20] (\QQ_in[21] [20]), 
            .\QQ_in[20][19] (\QQ_in[20] [19]), .\QQ_in[19][18] (\QQ_in[19] [18]), 
            .\QQ_in[18][17] (\QQ_in[18] [17]), .\QQ_in[17][16] (\QQ_in[17] [16]), 
            .\QQ_in[16][15] (\QQ_in[16] [15]), .\QQ_in[15][14] (\QQ_in[15] [14]), 
            .\QQ_in[14][13] (\QQ_in[14] [13]), .\QQ_in[13][12] (\QQ_in[13] [12]), 
            .\QQ_in[12][11] (\QQ_in[12] [11]), .\QQ_in[11][10] (\QQ_in[11] [10]), 
            .\QQ_in[10][9] (\QQ_in[10] [9]), .\QQ_in[9][8] (\QQ_in[9] [8]), 
            .\QQ_in[8][7] (\QQ_in[8] [7]), .\QQ_in[7][6] (\QQ_in[7] [6]), 
            .\QQ_in[6][5] (\QQ_in[6] [5]), .\QQ_in[24][23] (\QQ_in[24] [23]), 
            .\QQ_in[5][4] (\QQ_in[5] [4]), .\QQ_in[4][3] (\QQ_in[4] [3]), 
            .\QQ_in[3][2] (\QQ_in[3] [2]), .\QQ_in[2][1] (\QQ_in[2] [1]), 
            .\QQ_in[23][22] (\QQ_in[23] [22]), .GND_net(GND_net), .\B_int[21] (B_int[21]), 
            .\B_int[22] (B_int[22]), .\B_int[19] (B_int[19]), .\B_int[20] (B_int[20]), 
            .\B_int[17] (B_int[17]), .\B_int[18] (B_int[18]), .\B_int[15] (B_int[15]), 
            .\B_int[16] (B_int[16]), .\B_int[13] (B_int[13]), .\B_int[14] (B_int[14]), 
            .\B_int[11] (B_int[11]), .\B_int[12] (B_int[12]), .\B_int[9] (B_int[9]), 
            .\B_int[10] (B_int[10]), .\B_int[7] (B_int[7]), .\B_int[8] (B_int[8]), 
            .\B_int[5] (B_int[5]), .\B_int[6] (B_int[6]), .\B_int[3] (B_int[3]), 
            .\B_int[4] (B_int[4]), .\B_int[1] (B_int[1]), .\B_int[2] (B_int[2]), 
            .\B_int[0] (B_int[0]), .\QQ_in[1][0] (\QQ_in[1] [0]), .n9256(n9256), 
            .\QQ_in[25][24] (\QQ_in[25] [24]), .\QQ_in[26][25] (\QQ_in[26] [25]), 
            .\A_int[21] (A_int[21]), .\A_int[22] (A_int[22]), .\A_int[19] (A_int[19]), 
            .\A_int[20] (A_int[20]), .\A_int[17] (A_int[17]), .\A_int[18] (A_int[18]), 
            .\A_int[15] (A_int[15]), .\A_int[16] (A_int[16]), .\A_int[13] (A_int[13]), 
            .\A_int[14] (A_int[14]), .\A_int[11] (A_int[11]), .\A_int[12] (A_int[12]), 
            .\A_int[9] (A_int[9]), .\A_int[10] (A_int[10]), .\A_int[7] (A_int[7]), 
            .\A_int[8] (A_int[8]), .\A_int[5] (A_int[5]), .\A_int[6] (A_int[6]), 
            .\A_int[3] (A_int[3]), .\A_int[4] (A_int[4]), .\A_int[1] (A_int[1]), 
            .\A_int[2] (A_int[2]), .\A_int[0] (A_int[0]));
    
endmodule
//
// Verilog Description of module \div_nr_wsticky(24,27) 
//

module \div_nr_wsticky(24,27)  (\QQ_in[22][21] , \QQ_in[21][20] , \QQ_in[20][19] , 
            \QQ_in[19][18] , \QQ_in[18][17] , \QQ_in[17][16] , \QQ_in[16][15] , 
            \QQ_in[15][14] , \QQ_in[14][13] , \QQ_in[13][12] , \QQ_in[12][11] , 
            \QQ_in[11][10] , \QQ_in[10][9] , \QQ_in[9][8] , \QQ_in[8][7] , 
            \QQ_in[7][6] , \QQ_in[6][5] , \QQ_in[24][23] , \QQ_in[5][4] , 
            \QQ_in[4][3] , \QQ_in[3][2] , \QQ_in[2][1] , \QQ_in[23][22] , 
            GND_net, \B_int[21] , \B_int[22] , \B_int[19] , \B_int[20] , 
            \B_int[17] , \B_int[18] , \B_int[15] , \B_int[16] , \B_int[13] , 
            \B_int[14] , \B_int[11] , \B_int[12] , \B_int[9] , \B_int[10] , 
            \B_int[7] , \B_int[8] , \B_int[5] , \B_int[6] , \B_int[3] , 
            \B_int[4] , \B_int[1] , \B_int[2] , \B_int[0] , \QQ_in[1][0] , 
            n9256, \QQ_in[25][24] , \QQ_in[26][25] , \A_int[21] , \A_int[22] , 
            \A_int[19] , \A_int[20] , \A_int[17] , \A_int[18] , \A_int[15] , 
            \A_int[16] , \A_int[13] , \A_int[14] , \A_int[11] , \A_int[12] , 
            \A_int[9] , \A_int[10] , \A_int[7] , \A_int[8] , \A_int[5] , 
            \A_int[6] , \A_int[3] , \A_int[4] , \A_int[1] , \A_int[2] , 
            \A_int[0] );
    output \QQ_in[22][21] ;
    output \QQ_in[21][20] ;
    output \QQ_in[20][19] ;
    output \QQ_in[19][18] ;
    output \QQ_in[18][17] ;
    output \QQ_in[17][16] ;
    output \QQ_in[16][15] ;
    output \QQ_in[15][14] ;
    output \QQ_in[14][13] ;
    output \QQ_in[13][12] ;
    output \QQ_in[12][11] ;
    output \QQ_in[11][10] ;
    output \QQ_in[10][9] ;
    output \QQ_in[9][8] ;
    output \QQ_in[8][7] ;
    output \QQ_in[7][6] ;
    output \QQ_in[6][5] ;
    output \QQ_in[24][23] ;
    output \QQ_in[5][4] ;
    output \QQ_in[4][3] ;
    output \QQ_in[3][2] ;
    output \QQ_in[2][1] ;
    output \QQ_in[23][22] ;
    input GND_net;
    input \B_int[21] ;
    input \B_int[22] ;
    input \B_int[19] ;
    input \B_int[20] ;
    input \B_int[17] ;
    input \B_int[18] ;
    input \B_int[15] ;
    input \B_int[16] ;
    input \B_int[13] ;
    input \B_int[14] ;
    input \B_int[11] ;
    input \B_int[12] ;
    input \B_int[9] ;
    input \B_int[10] ;
    input \B_int[7] ;
    input \B_int[8] ;
    input \B_int[5] ;
    input \B_int[6] ;
    input \B_int[3] ;
    input \B_int[4] ;
    input \B_int[1] ;
    input \B_int[2] ;
    input \B_int[0] ;
    output \QQ_in[1][0] ;
    input n9256;
    output \QQ_in[25][24] ;
    output \QQ_in[26][25] ;
    input \A_int[21] ;
    input \A_int[22] ;
    input \A_int[19] ;
    input \A_int[20] ;
    input \A_int[17] ;
    input \A_int[18] ;
    input \A_int[15] ;
    input \A_int[16] ;
    input \A_int[13] ;
    input \A_int[14] ;
    input \A_int[11] ;
    input \A_int[12] ;
    input \A_int[9] ;
    input \A_int[10] ;
    input \A_int[7] ;
    input \A_int[8] ;
    input \A_int[5] ;
    input \A_int[6] ;
    input \A_int[3] ;
    input \A_int[4] ;
    input \A_int[1] ;
    input \A_int[2] ;
    input \A_int[0] ;
    
    wire [26:0]frac_div;   // c:/users/yisong/documents/new/mlp/fp_div.vhd(72[11:19])
    wire [24:0]\m_cablesIn[8] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[9] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[7] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[6] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[5] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[4] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[3] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[2] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[1] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[25] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[24] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[23] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[22] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[21] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[20] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[19] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[18] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[17] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[16] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[15] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[14] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[13] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[12] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[11] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    wire [24:0]\m_cablesIn[10] ;   // c:/users/yisong/documents/new/mlp/div_nr_wsticky.vhd(45[11:21])
    
    LUT4 i9_1_lut (.A(\QQ_in[22][21] ), .Z(frac_div[5])) /* synthesis lut_function=(!(A)) */ ;
    defparam i9_1_lut.init = 16'h5555;
    LUT4 i10_1_lut (.A(\QQ_in[21][20] ), .Z(frac_div[6])) /* synthesis lut_function=(!(A)) */ ;
    defparam i10_1_lut.init = 16'h5555;
    LUT4 i11_1_lut (.A(\QQ_in[20][19] ), .Z(frac_div[7])) /* synthesis lut_function=(!(A)) */ ;
    defparam i11_1_lut.init = 16'h5555;
    LUT4 i12_1_lut (.A(\QQ_in[19][18] ), .Z(frac_div[8])) /* synthesis lut_function=(!(A)) */ ;
    defparam i12_1_lut.init = 16'h5555;
    LUT4 i13_1_lut (.A(\QQ_in[18][17] ), .Z(frac_div[9])) /* synthesis lut_function=(!(A)) */ ;
    defparam i13_1_lut.init = 16'h5555;
    LUT4 i14_1_lut (.A(\QQ_in[17][16] ), .Z(frac_div[10])) /* synthesis lut_function=(!(A)) */ ;
    defparam i14_1_lut.init = 16'h5555;
    LUT4 i15_1_lut (.A(\QQ_in[16][15] ), .Z(frac_div[11])) /* synthesis lut_function=(!(A)) */ ;
    defparam i15_1_lut.init = 16'h5555;
    LUT4 i16_1_lut (.A(\QQ_in[15][14] ), .Z(frac_div[12])) /* synthesis lut_function=(!(A)) */ ;
    defparam i16_1_lut.init = 16'h5555;
    LUT4 i17_1_lut (.A(\QQ_in[14][13] ), .Z(frac_div[13])) /* synthesis lut_function=(!(A)) */ ;
    defparam i17_1_lut.init = 16'h5555;
    LUT4 i18_1_lut (.A(\QQ_in[13][12] ), .Z(frac_div[14])) /* synthesis lut_function=(!(A)) */ ;
    defparam i18_1_lut.init = 16'h5555;
    LUT4 i19_1_lut (.A(\QQ_in[12][11] ), .Z(frac_div[15])) /* synthesis lut_function=(!(A)) */ ;
    defparam i19_1_lut.init = 16'h5555;
    LUT4 i20_1_lut (.A(\QQ_in[11][10] ), .Z(frac_div[16])) /* synthesis lut_function=(!(A)) */ ;
    defparam i20_1_lut.init = 16'h5555;
    LUT4 i21_1_lut (.A(\QQ_in[10][9] ), .Z(frac_div[17])) /* synthesis lut_function=(!(A)) */ ;
    defparam i21_1_lut.init = 16'h5555;
    LUT4 i22_1_lut (.A(\QQ_in[9][8] ), .Z(frac_div[18])) /* synthesis lut_function=(!(A)) */ ;
    defparam i22_1_lut.init = 16'h5555;
    LUT4 i23_1_lut (.A(\QQ_in[8][7] ), .Z(frac_div[19])) /* synthesis lut_function=(!(A)) */ ;
    defparam i23_1_lut.init = 16'h5555;
    LUT4 i24_1_lut (.A(\QQ_in[7][6] ), .Z(frac_div[20])) /* synthesis lut_function=(!(A)) */ ;
    defparam i24_1_lut.init = 16'h5555;
    LUT4 i25_1_lut (.A(\QQ_in[6][5] ), .Z(frac_div[21])) /* synthesis lut_function=(!(A)) */ ;
    defparam i25_1_lut.init = 16'h5555;
    LUT4 i7_1_lut (.A(\QQ_in[24][23] ), .Z(frac_div[3])) /* synthesis lut_function=(!(A)) */ ;
    defparam i7_1_lut.init = 16'h5555;
    LUT4 i26_1_lut (.A(\QQ_in[5][4] ), .Z(frac_div[22])) /* synthesis lut_function=(!(A)) */ ;
    defparam i26_1_lut.init = 16'h5555;
    LUT4 i27_1_lut (.A(\QQ_in[4][3] ), .Z(frac_div[23])) /* synthesis lut_function=(!(A)) */ ;
    defparam i27_1_lut.init = 16'h5555;
    LUT4 i28_1_lut (.A(\QQ_in[3][2] ), .Z(frac_div[24])) /* synthesis lut_function=(!(A)) */ ;
    defparam i28_1_lut.init = 16'h5555;
    LUT4 i29_1_lut (.A(\QQ_in[2][1] ), .Z(frac_div[25])) /* synthesis lut_function=(!(A)) */ ;
    defparam i29_1_lut.init = 16'h5555;
    LUT4 i8_1_lut (.A(\QQ_in[23][22] ), .Z(frac_div[4])) /* synthesis lut_function=(!(A)) */ ;
    defparam i8_1_lut.init = 16'h5555;
    \a_s(24)  \divisor_9..int_mod  (.\m_cablesIn[8][23] (\m_cablesIn[8] [23]), 
            .\QQ_in[8][7] (\QQ_in[8][7] ), .GND_net(GND_net), .\m_cablesIn[8][24] (\m_cablesIn[8] [24]), 
            .\m_cablesIn[9][24] (\m_cablesIn[9] [24]), .\QQ_in[9][8] (\QQ_in[9][8] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[8][21] (\m_cablesIn[8] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[8][22] (\m_cablesIn[8] [22]), 
            .\m_cablesIn[9][22] (\m_cablesIn[9] [22]), .\m_cablesIn[9][23] (\m_cablesIn[9] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[8][19] (\m_cablesIn[8] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[8][20] (\m_cablesIn[8] [20]), 
            .\m_cablesIn[9][20] (\m_cablesIn[9] [20]), .\m_cablesIn[9][21] (\m_cablesIn[9] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[8][17] (\m_cablesIn[8] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[8][18] (\m_cablesIn[8] [18]), 
            .\m_cablesIn[9][18] (\m_cablesIn[9] [18]), .\m_cablesIn[9][19] (\m_cablesIn[9] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[8][15] (\m_cablesIn[8] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[8][16] (\m_cablesIn[8] [16]), 
            .\m_cablesIn[9][16] (\m_cablesIn[9] [16]), .\m_cablesIn[9][17] (\m_cablesIn[9] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[8][13] (\m_cablesIn[8] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[8][14] (\m_cablesIn[8] [14]), 
            .\m_cablesIn[9][14] (\m_cablesIn[9] [14]), .\m_cablesIn[9][15] (\m_cablesIn[9] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[8][11] (\m_cablesIn[8] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[8][12] (\m_cablesIn[8] [12]), 
            .\m_cablesIn[9][12] (\m_cablesIn[9] [12]), .\m_cablesIn[9][13] (\m_cablesIn[9] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[8][9] (\m_cablesIn[8] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[8][10] (\m_cablesIn[8] [10]), 
            .\m_cablesIn[9][10] (\m_cablesIn[9] [10]), .\m_cablesIn[9][11] (\m_cablesIn[9] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[8][7] (\m_cablesIn[8] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[8][8] (\m_cablesIn[8] [8]), 
            .\m_cablesIn[9][8] (\m_cablesIn[9] [8]), .\m_cablesIn[9][9] (\m_cablesIn[9] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[8][5] (\m_cablesIn[8] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[8][6] (\m_cablesIn[8] [6]), 
            .\m_cablesIn[9][6] (\m_cablesIn[9] [6]), .\m_cablesIn[9][7] (\m_cablesIn[9] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[8][3] (\m_cablesIn[8] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[8][4] (\m_cablesIn[8] [4]), 
            .\m_cablesIn[9][4] (\m_cablesIn[9] [4]), .\m_cablesIn[9][5] (\m_cablesIn[9] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[8][1] (\m_cablesIn[8] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[8][2] (\m_cablesIn[8] [2]), 
            .\m_cablesIn[9][2] (\m_cablesIn[9] [2]), .\m_cablesIn[9][3] (\m_cablesIn[9] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[19] (frac_div[19]), .\m_cablesIn[9][1] (\m_cablesIn[9] [1]));
    \a_s(24)_U0  \divisor_8..int_mod  (.\m_cablesIn[7][23] (\m_cablesIn[7] [23]), 
            .\QQ_in[7][6] (\QQ_in[7][6] ), .GND_net(GND_net), .\m_cablesIn[7][24] (\m_cablesIn[7] [24]), 
            .\m_cablesIn[8][24] (\m_cablesIn[8] [24]), .\QQ_in[8][7] (\QQ_in[8][7] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[7][21] (\m_cablesIn[7] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[7][22] (\m_cablesIn[7] [22]), 
            .\m_cablesIn[8][22] (\m_cablesIn[8] [22]), .\m_cablesIn[8][23] (\m_cablesIn[8] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[7][19] (\m_cablesIn[7] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[7][20] (\m_cablesIn[7] [20]), 
            .\m_cablesIn[8][20] (\m_cablesIn[8] [20]), .\m_cablesIn[8][21] (\m_cablesIn[8] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[7][17] (\m_cablesIn[7] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[7][18] (\m_cablesIn[7] [18]), 
            .\m_cablesIn[8][18] (\m_cablesIn[8] [18]), .\m_cablesIn[8][19] (\m_cablesIn[8] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[7][15] (\m_cablesIn[7] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[7][16] (\m_cablesIn[7] [16]), 
            .\m_cablesIn[8][16] (\m_cablesIn[8] [16]), .\m_cablesIn[8][17] (\m_cablesIn[8] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[7][13] (\m_cablesIn[7] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[7][14] (\m_cablesIn[7] [14]), 
            .\m_cablesIn[8][14] (\m_cablesIn[8] [14]), .\m_cablesIn[8][15] (\m_cablesIn[8] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[7][11] (\m_cablesIn[7] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[7][12] (\m_cablesIn[7] [12]), 
            .\m_cablesIn[8][12] (\m_cablesIn[8] [12]), .\m_cablesIn[8][13] (\m_cablesIn[8] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[7][9] (\m_cablesIn[7] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[7][10] (\m_cablesIn[7] [10]), 
            .\m_cablesIn[8][10] (\m_cablesIn[8] [10]), .\m_cablesIn[8][11] (\m_cablesIn[8] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[7][7] (\m_cablesIn[7] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[7][8] (\m_cablesIn[7] [8]), 
            .\m_cablesIn[8][8] (\m_cablesIn[8] [8]), .\m_cablesIn[8][9] (\m_cablesIn[8] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[7][5] (\m_cablesIn[7] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[7][6] (\m_cablesIn[7] [6]), 
            .\m_cablesIn[8][6] (\m_cablesIn[8] [6]), .\m_cablesIn[8][7] (\m_cablesIn[8] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[7][3] (\m_cablesIn[7] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[7][4] (\m_cablesIn[7] [4]), 
            .\m_cablesIn[8][4] (\m_cablesIn[8] [4]), .\m_cablesIn[8][5] (\m_cablesIn[8] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[7][1] (\m_cablesIn[7] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[7][2] (\m_cablesIn[7] [2]), 
            .\m_cablesIn[8][2] (\m_cablesIn[8] [2]), .\m_cablesIn[8][3] (\m_cablesIn[8] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[20] (frac_div[20]), .\m_cablesIn[8][1] (\m_cablesIn[8] [1]));
    \a_s(24)_U1  \divisor_7..int_mod  (.\m_cablesIn[6][23] (\m_cablesIn[6] [23]), 
            .\QQ_in[6][5] (\QQ_in[6][5] ), .GND_net(GND_net), .\m_cablesIn[6][24] (\m_cablesIn[6] [24]), 
            .\m_cablesIn[7][24] (\m_cablesIn[7] [24]), .\QQ_in[7][6] (\QQ_in[7][6] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[6][21] (\m_cablesIn[6] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[6][22] (\m_cablesIn[6] [22]), 
            .\m_cablesIn[7][22] (\m_cablesIn[7] [22]), .\m_cablesIn[7][23] (\m_cablesIn[7] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[6][19] (\m_cablesIn[6] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[6][20] (\m_cablesIn[6] [20]), 
            .\m_cablesIn[7][20] (\m_cablesIn[7] [20]), .\m_cablesIn[7][21] (\m_cablesIn[7] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[6][17] (\m_cablesIn[6] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[6][18] (\m_cablesIn[6] [18]), 
            .\m_cablesIn[7][18] (\m_cablesIn[7] [18]), .\m_cablesIn[7][19] (\m_cablesIn[7] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[6][15] (\m_cablesIn[6] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[6][16] (\m_cablesIn[6] [16]), 
            .\m_cablesIn[7][16] (\m_cablesIn[7] [16]), .\m_cablesIn[7][17] (\m_cablesIn[7] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[6][13] (\m_cablesIn[6] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[6][14] (\m_cablesIn[6] [14]), 
            .\m_cablesIn[7][14] (\m_cablesIn[7] [14]), .\m_cablesIn[7][15] (\m_cablesIn[7] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[6][11] (\m_cablesIn[6] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[6][12] (\m_cablesIn[6] [12]), 
            .\m_cablesIn[7][12] (\m_cablesIn[7] [12]), .\m_cablesIn[7][13] (\m_cablesIn[7] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[6][9] (\m_cablesIn[6] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[6][10] (\m_cablesIn[6] [10]), 
            .\m_cablesIn[7][10] (\m_cablesIn[7] [10]), .\m_cablesIn[7][11] (\m_cablesIn[7] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[6][7] (\m_cablesIn[6] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[6][8] (\m_cablesIn[6] [8]), 
            .\m_cablesIn[7][8] (\m_cablesIn[7] [8]), .\m_cablesIn[7][9] (\m_cablesIn[7] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[6][5] (\m_cablesIn[6] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[6][6] (\m_cablesIn[6] [6]), 
            .\m_cablesIn[7][6] (\m_cablesIn[7] [6]), .\m_cablesIn[7][7] (\m_cablesIn[7] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[6][3] (\m_cablesIn[6] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[6][4] (\m_cablesIn[6] [4]), 
            .\m_cablesIn[7][4] (\m_cablesIn[7] [4]), .\m_cablesIn[7][5] (\m_cablesIn[7] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[6][1] (\m_cablesIn[6] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[6][2] (\m_cablesIn[6] [2]), 
            .\m_cablesIn[7][2] (\m_cablesIn[7] [2]), .\m_cablesIn[7][3] (\m_cablesIn[7] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[21] (frac_div[21]), .\m_cablesIn[7][1] (\m_cablesIn[7] [1]));
    \a_s(24)_U2  \divisor_6..int_mod  (.\m_cablesIn[5][23] (\m_cablesIn[5] [23]), 
            .\QQ_in[5][4] (\QQ_in[5][4] ), .GND_net(GND_net), .\m_cablesIn[5][24] (\m_cablesIn[5] [24]), 
            .\m_cablesIn[6][24] (\m_cablesIn[6] [24]), .\QQ_in[6][5] (\QQ_in[6][5] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[5][21] (\m_cablesIn[5] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[5][22] (\m_cablesIn[5] [22]), 
            .\m_cablesIn[6][22] (\m_cablesIn[6] [22]), .\m_cablesIn[6][23] (\m_cablesIn[6] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[5][19] (\m_cablesIn[5] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[5][20] (\m_cablesIn[5] [20]), 
            .\m_cablesIn[6][20] (\m_cablesIn[6] [20]), .\m_cablesIn[6][21] (\m_cablesIn[6] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[5][17] (\m_cablesIn[5] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[5][18] (\m_cablesIn[5] [18]), 
            .\m_cablesIn[6][18] (\m_cablesIn[6] [18]), .\m_cablesIn[6][19] (\m_cablesIn[6] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[5][15] (\m_cablesIn[5] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[5][16] (\m_cablesIn[5] [16]), 
            .\m_cablesIn[6][16] (\m_cablesIn[6] [16]), .\m_cablesIn[6][17] (\m_cablesIn[6] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[5][13] (\m_cablesIn[5] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[5][14] (\m_cablesIn[5] [14]), 
            .\m_cablesIn[6][14] (\m_cablesIn[6] [14]), .\m_cablesIn[6][15] (\m_cablesIn[6] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[5][11] (\m_cablesIn[5] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[5][12] (\m_cablesIn[5] [12]), 
            .\m_cablesIn[6][12] (\m_cablesIn[6] [12]), .\m_cablesIn[6][13] (\m_cablesIn[6] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[5][9] (\m_cablesIn[5] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[5][10] (\m_cablesIn[5] [10]), 
            .\m_cablesIn[6][10] (\m_cablesIn[6] [10]), .\m_cablesIn[6][11] (\m_cablesIn[6] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[5][7] (\m_cablesIn[5] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[5][8] (\m_cablesIn[5] [8]), 
            .\m_cablesIn[6][8] (\m_cablesIn[6] [8]), .\m_cablesIn[6][9] (\m_cablesIn[6] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[5][5] (\m_cablesIn[5] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[5][6] (\m_cablesIn[5] [6]), 
            .\m_cablesIn[6][6] (\m_cablesIn[6] [6]), .\m_cablesIn[6][7] (\m_cablesIn[6] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[5][3] (\m_cablesIn[5] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[5][4] (\m_cablesIn[5] [4]), 
            .\m_cablesIn[6][4] (\m_cablesIn[6] [4]), .\m_cablesIn[6][5] (\m_cablesIn[6] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[5][1] (\m_cablesIn[5] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[5][2] (\m_cablesIn[5] [2]), 
            .\m_cablesIn[6][2] (\m_cablesIn[6] [2]), .\m_cablesIn[6][3] (\m_cablesIn[6] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[22] (frac_div[22]), .\m_cablesIn[6][1] (\m_cablesIn[6] [1]));
    \a_s(24)_U3  \divisor_5..int_mod  (.\m_cablesIn[4][23] (\m_cablesIn[4] [23]), 
            .\QQ_in[4][3] (\QQ_in[4][3] ), .GND_net(GND_net), .\m_cablesIn[4][24] (\m_cablesIn[4] [24]), 
            .\m_cablesIn[5][24] (\m_cablesIn[5] [24]), .\QQ_in[5][4] (\QQ_in[5][4] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[4][21] (\m_cablesIn[4] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[4][22] (\m_cablesIn[4] [22]), 
            .\m_cablesIn[5][22] (\m_cablesIn[5] [22]), .\m_cablesIn[5][23] (\m_cablesIn[5] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[4][19] (\m_cablesIn[4] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[4][20] (\m_cablesIn[4] [20]), 
            .\m_cablesIn[5][20] (\m_cablesIn[5] [20]), .\m_cablesIn[5][21] (\m_cablesIn[5] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[4][17] (\m_cablesIn[4] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[4][18] (\m_cablesIn[4] [18]), 
            .\m_cablesIn[5][18] (\m_cablesIn[5] [18]), .\m_cablesIn[5][19] (\m_cablesIn[5] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[4][15] (\m_cablesIn[4] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[4][16] (\m_cablesIn[4] [16]), 
            .\m_cablesIn[5][16] (\m_cablesIn[5] [16]), .\m_cablesIn[5][17] (\m_cablesIn[5] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[4][13] (\m_cablesIn[4] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[4][14] (\m_cablesIn[4] [14]), 
            .\m_cablesIn[5][14] (\m_cablesIn[5] [14]), .\m_cablesIn[5][15] (\m_cablesIn[5] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[4][11] (\m_cablesIn[4] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[4][12] (\m_cablesIn[4] [12]), 
            .\m_cablesIn[5][12] (\m_cablesIn[5] [12]), .\m_cablesIn[5][13] (\m_cablesIn[5] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[4][9] (\m_cablesIn[4] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[4][10] (\m_cablesIn[4] [10]), 
            .\m_cablesIn[5][10] (\m_cablesIn[5] [10]), .\m_cablesIn[5][11] (\m_cablesIn[5] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[4][7] (\m_cablesIn[4] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[4][8] (\m_cablesIn[4] [8]), 
            .\m_cablesIn[5][8] (\m_cablesIn[5] [8]), .\m_cablesIn[5][9] (\m_cablesIn[5] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[4][5] (\m_cablesIn[4] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[4][6] (\m_cablesIn[4] [6]), 
            .\m_cablesIn[5][6] (\m_cablesIn[5] [6]), .\m_cablesIn[5][7] (\m_cablesIn[5] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[4][3] (\m_cablesIn[4] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[4][4] (\m_cablesIn[4] [4]), 
            .\m_cablesIn[5][4] (\m_cablesIn[5] [4]), .\m_cablesIn[5][5] (\m_cablesIn[5] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[4][1] (\m_cablesIn[4] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[4][2] (\m_cablesIn[4] [2]), 
            .\m_cablesIn[5][2] (\m_cablesIn[5] [2]), .\m_cablesIn[5][3] (\m_cablesIn[5] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[23] (frac_div[23]), .\m_cablesIn[5][1] (\m_cablesIn[5] [1]));
    \a_s(24)_U4  \divisor_4..int_mod  (.\m_cablesIn[3][23] (\m_cablesIn[3] [23]), 
            .\QQ_in[3][2] (\QQ_in[3][2] ), .GND_net(GND_net), .\m_cablesIn[3][24] (\m_cablesIn[3] [24]), 
            .\m_cablesIn[4][24] (\m_cablesIn[4] [24]), .\QQ_in[4][3] (\QQ_in[4][3] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[3][21] (\m_cablesIn[3] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[3][22] (\m_cablesIn[3] [22]), 
            .\m_cablesIn[4][22] (\m_cablesIn[4] [22]), .\m_cablesIn[4][23] (\m_cablesIn[4] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[3][19] (\m_cablesIn[3] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[3][20] (\m_cablesIn[3] [20]), 
            .\m_cablesIn[4][20] (\m_cablesIn[4] [20]), .\m_cablesIn[4][21] (\m_cablesIn[4] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[3][17] (\m_cablesIn[3] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[3][18] (\m_cablesIn[3] [18]), 
            .\m_cablesIn[4][18] (\m_cablesIn[4] [18]), .\m_cablesIn[4][19] (\m_cablesIn[4] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[3][15] (\m_cablesIn[3] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[3][16] (\m_cablesIn[3] [16]), 
            .\m_cablesIn[4][16] (\m_cablesIn[4] [16]), .\m_cablesIn[4][17] (\m_cablesIn[4] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[3][13] (\m_cablesIn[3] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[3][14] (\m_cablesIn[3] [14]), 
            .\m_cablesIn[4][14] (\m_cablesIn[4] [14]), .\m_cablesIn[4][15] (\m_cablesIn[4] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[3][11] (\m_cablesIn[3] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[3][12] (\m_cablesIn[3] [12]), 
            .\m_cablesIn[4][12] (\m_cablesIn[4] [12]), .\m_cablesIn[4][13] (\m_cablesIn[4] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[3][9] (\m_cablesIn[3] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[3][10] (\m_cablesIn[3] [10]), 
            .\m_cablesIn[4][10] (\m_cablesIn[4] [10]), .\m_cablesIn[4][11] (\m_cablesIn[4] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[3][7] (\m_cablesIn[3] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[3][8] (\m_cablesIn[3] [8]), 
            .\m_cablesIn[4][8] (\m_cablesIn[4] [8]), .\m_cablesIn[4][9] (\m_cablesIn[4] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[3][5] (\m_cablesIn[3] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[3][6] (\m_cablesIn[3] [6]), 
            .\m_cablesIn[4][6] (\m_cablesIn[4] [6]), .\m_cablesIn[4][7] (\m_cablesIn[4] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[3][3] (\m_cablesIn[3] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[3][4] (\m_cablesIn[3] [4]), 
            .\m_cablesIn[4][4] (\m_cablesIn[4] [4]), .\m_cablesIn[4][5] (\m_cablesIn[4] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[3][1] (\m_cablesIn[3] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[3][2] (\m_cablesIn[3] [2]), 
            .\m_cablesIn[4][2] (\m_cablesIn[4] [2]), .\m_cablesIn[4][3] (\m_cablesIn[4] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[24] (frac_div[24]), .\m_cablesIn[4][1] (\m_cablesIn[4] [1]));
    \a_s(24)_U5  \divisor_3..int_mod  (.\m_cablesIn[2][23] (\m_cablesIn[2] [23]), 
            .\QQ_in[2][1] (\QQ_in[2][1] ), .GND_net(GND_net), .\m_cablesIn[2][24] (\m_cablesIn[2] [24]), 
            .\m_cablesIn[3][24] (\m_cablesIn[3] [24]), .\QQ_in[3][2] (\QQ_in[3][2] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[2][21] (\m_cablesIn[2] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[2][22] (\m_cablesIn[2] [22]), 
            .\m_cablesIn[3][22] (\m_cablesIn[3] [22]), .\m_cablesIn[3][23] (\m_cablesIn[3] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[2][19] (\m_cablesIn[2] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[2][20] (\m_cablesIn[2] [20]), 
            .\m_cablesIn[3][20] (\m_cablesIn[3] [20]), .\m_cablesIn[3][21] (\m_cablesIn[3] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[2][17] (\m_cablesIn[2] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[2][18] (\m_cablesIn[2] [18]), 
            .\m_cablesIn[3][18] (\m_cablesIn[3] [18]), .\m_cablesIn[3][19] (\m_cablesIn[3] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[2][15] (\m_cablesIn[2] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[2][16] (\m_cablesIn[2] [16]), 
            .\m_cablesIn[3][16] (\m_cablesIn[3] [16]), .\m_cablesIn[3][17] (\m_cablesIn[3] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[2][13] (\m_cablesIn[2] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[2][14] (\m_cablesIn[2] [14]), 
            .\m_cablesIn[3][14] (\m_cablesIn[3] [14]), .\m_cablesIn[3][15] (\m_cablesIn[3] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[2][11] (\m_cablesIn[2] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[2][12] (\m_cablesIn[2] [12]), 
            .\m_cablesIn[3][12] (\m_cablesIn[3] [12]), .\m_cablesIn[3][13] (\m_cablesIn[3] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[2][9] (\m_cablesIn[2] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[2][10] (\m_cablesIn[2] [10]), 
            .\m_cablesIn[3][10] (\m_cablesIn[3] [10]), .\m_cablesIn[3][11] (\m_cablesIn[3] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[2][7] (\m_cablesIn[2] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[2][8] (\m_cablesIn[2] [8]), 
            .\m_cablesIn[3][8] (\m_cablesIn[3] [8]), .\m_cablesIn[3][9] (\m_cablesIn[3] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[2][5] (\m_cablesIn[2] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[2][6] (\m_cablesIn[2] [6]), 
            .\m_cablesIn[3][6] (\m_cablesIn[3] [6]), .\m_cablesIn[3][7] (\m_cablesIn[3] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[2][3] (\m_cablesIn[2] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[2][4] (\m_cablesIn[2] [4]), 
            .\m_cablesIn[3][4] (\m_cablesIn[3] [4]), .\m_cablesIn[3][5] (\m_cablesIn[3] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[2][1] (\m_cablesIn[2] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[2][2] (\m_cablesIn[2] [2]), 
            .\m_cablesIn[3][2] (\m_cablesIn[3] [2]), .\m_cablesIn[3][3] (\m_cablesIn[3] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[25] (frac_div[25]), .\m_cablesIn[3][1] (\m_cablesIn[3] [1]));
    \a_s(24)_U6  \divisor_2..int_mod  (.\m_cablesIn[1][23] (\m_cablesIn[1] [23]), 
            .\QQ_in[1][0] (\QQ_in[1][0] ), .GND_net(GND_net), .\m_cablesIn[1][24] (\m_cablesIn[1] [24]), 
            .\m_cablesIn[2][24] (\m_cablesIn[2] [24]), .\QQ_in[2][1] (\QQ_in[2][1] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[1][21] (\m_cablesIn[1] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[1][22] (\m_cablesIn[1] [22]), 
            .\m_cablesIn[2][22] (\m_cablesIn[2] [22]), .\m_cablesIn[2][23] (\m_cablesIn[2] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[1][19] (\m_cablesIn[1] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[1][20] (\m_cablesIn[1] [20]), 
            .\m_cablesIn[2][20] (\m_cablesIn[2] [20]), .\m_cablesIn[2][21] (\m_cablesIn[2] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[1][17] (\m_cablesIn[1] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[1][18] (\m_cablesIn[1] [18]), 
            .\m_cablesIn[2][18] (\m_cablesIn[2] [18]), .\m_cablesIn[2][19] (\m_cablesIn[2] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[1][15] (\m_cablesIn[1] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[1][16] (\m_cablesIn[1] [16]), 
            .\m_cablesIn[2][16] (\m_cablesIn[2] [16]), .\m_cablesIn[2][17] (\m_cablesIn[2] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[1][13] (\m_cablesIn[1] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[1][14] (\m_cablesIn[1] [14]), 
            .\m_cablesIn[2][14] (\m_cablesIn[2] [14]), .\m_cablesIn[2][15] (\m_cablesIn[2] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[1][11] (\m_cablesIn[1] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[1][12] (\m_cablesIn[1] [12]), 
            .\m_cablesIn[2][12] (\m_cablesIn[2] [12]), .\m_cablesIn[2][13] (\m_cablesIn[2] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[1][9] (\m_cablesIn[1] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[1][10] (\m_cablesIn[1] [10]), 
            .\m_cablesIn[2][10] (\m_cablesIn[2] [10]), .\m_cablesIn[2][11] (\m_cablesIn[2] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[1][7] (\m_cablesIn[1] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[1][8] (\m_cablesIn[1] [8]), 
            .\m_cablesIn[2][8] (\m_cablesIn[2] [8]), .\m_cablesIn[2][9] (\m_cablesIn[2] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[1][5] (\m_cablesIn[1] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[1][6] (\m_cablesIn[1] [6]), 
            .\m_cablesIn[2][6] (\m_cablesIn[2] [6]), .\m_cablesIn[2][7] (\m_cablesIn[2] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[1][3] (\m_cablesIn[1] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[1][4] (\m_cablesIn[1] [4]), 
            .\m_cablesIn[2][4] (\m_cablesIn[2] [4]), .\m_cablesIn[2][5] (\m_cablesIn[2] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[1][1] (\m_cablesIn[1] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[1][2] (\m_cablesIn[1] [2]), 
            .\m_cablesIn[2][2] (\m_cablesIn[2] [2]), .\m_cablesIn[2][3] (\m_cablesIn[2] [3]), 
            .\B_int[0] (\B_int[0] ), .n9256(n9256), .\m_cablesIn[2][1] (\m_cablesIn[2] [1]));
    \a_s(24)_U7  \divisor_26..int_mod  (.\m_cablesIn[25][23] (\m_cablesIn[25] [23]), 
            .\QQ_in[25][24] (\QQ_in[25][24] ), .GND_net(GND_net), .\m_cablesIn[25][24] (\m_cablesIn[25] [24]), 
            .\QQ_in[26][25] (\QQ_in[26][25] ), .\B_int[21] (\B_int[21] ), 
            .\m_cablesIn[25][21] (\m_cablesIn[25] [21]), .\B_int[22] (\B_int[22] ), 
            .\m_cablesIn[25][22] (\m_cablesIn[25] [22]), .\B_int[19] (\B_int[19] ), 
            .\m_cablesIn[25][19] (\m_cablesIn[25] [19]), .\B_int[20] (\B_int[20] ), 
            .\m_cablesIn[25][20] (\m_cablesIn[25] [20]), .\B_int[17] (\B_int[17] ), 
            .\m_cablesIn[25][17] (\m_cablesIn[25] [17]), .\B_int[18] (\B_int[18] ), 
            .\m_cablesIn[25][18] (\m_cablesIn[25] [18]), .\B_int[15] (\B_int[15] ), 
            .\m_cablesIn[25][15] (\m_cablesIn[25] [15]), .\B_int[16] (\B_int[16] ), 
            .\m_cablesIn[25][16] (\m_cablesIn[25] [16]), .\B_int[13] (\B_int[13] ), 
            .\m_cablesIn[25][13] (\m_cablesIn[25] [13]), .\B_int[14] (\B_int[14] ), 
            .\m_cablesIn[25][14] (\m_cablesIn[25] [14]), .\B_int[11] (\B_int[11] ), 
            .\m_cablesIn[25][11] (\m_cablesIn[25] [11]), .\B_int[12] (\B_int[12] ), 
            .\m_cablesIn[25][12] (\m_cablesIn[25] [12]), .\B_int[9] (\B_int[9] ), 
            .\m_cablesIn[25][9] (\m_cablesIn[25] [9]), .\B_int[10] (\B_int[10] ), 
            .\m_cablesIn[25][10] (\m_cablesIn[25] [10]), .\B_int[7] (\B_int[7] ), 
            .\m_cablesIn[25][7] (\m_cablesIn[25] [7]), .\B_int[8] (\B_int[8] ), 
            .\m_cablesIn[25][8] (\m_cablesIn[25] [8]), .\B_int[5] (\B_int[5] ), 
            .\m_cablesIn[25][5] (\m_cablesIn[25] [5]), .\B_int[6] (\B_int[6] ), 
            .\m_cablesIn[25][6] (\m_cablesIn[25] [6]), .\B_int[3] (\B_int[3] ), 
            .\m_cablesIn[25][3] (\m_cablesIn[25] [3]), .\B_int[4] (\B_int[4] ), 
            .\m_cablesIn[25][4] (\m_cablesIn[25] [4]), .\B_int[1] (\B_int[1] ), 
            .\m_cablesIn[25][1] (\m_cablesIn[25] [1]), .\B_int[2] (\B_int[2] ), 
            .\m_cablesIn[25][2] (\m_cablesIn[25] [2]), .\B_int[0] (\B_int[0] ), 
            .\frac_div[2] (frac_div[2]));
    \a_s(24)_U8  \divisor_25..int_mod  (.\QQ_in[25][24] (\QQ_in[25][24] ), 
            .\frac_div[2] (frac_div[2]), .\m_cablesIn[24][23] (\m_cablesIn[24] [23]), 
            .\QQ_in[24][23] (\QQ_in[24][23] ), .GND_net(GND_net), .\m_cablesIn[24][24] (\m_cablesIn[24] [24]), 
            .\m_cablesIn[25][24] (\m_cablesIn[25] [24]), .\B_int[21] (\B_int[21] ), 
            .\m_cablesIn[24][21] (\m_cablesIn[24] [21]), .\B_int[22] (\B_int[22] ), 
            .\m_cablesIn[24][22] (\m_cablesIn[24] [22]), .\m_cablesIn[25][22] (\m_cablesIn[25] [22]), 
            .\m_cablesIn[25][23] (\m_cablesIn[25] [23]), .\B_int[19] (\B_int[19] ), 
            .\m_cablesIn[24][19] (\m_cablesIn[24] [19]), .\B_int[20] (\B_int[20] ), 
            .\m_cablesIn[24][20] (\m_cablesIn[24] [20]), .\m_cablesIn[25][20] (\m_cablesIn[25] [20]), 
            .\m_cablesIn[25][21] (\m_cablesIn[25] [21]), .\B_int[17] (\B_int[17] ), 
            .\m_cablesIn[24][17] (\m_cablesIn[24] [17]), .\B_int[18] (\B_int[18] ), 
            .\m_cablesIn[24][18] (\m_cablesIn[24] [18]), .\m_cablesIn[25][18] (\m_cablesIn[25] [18]), 
            .\m_cablesIn[25][19] (\m_cablesIn[25] [19]), .\B_int[15] (\B_int[15] ), 
            .\m_cablesIn[24][15] (\m_cablesIn[24] [15]), .\B_int[16] (\B_int[16] ), 
            .\m_cablesIn[24][16] (\m_cablesIn[24] [16]), .\m_cablesIn[25][16] (\m_cablesIn[25] [16]), 
            .\m_cablesIn[25][17] (\m_cablesIn[25] [17]), .\B_int[13] (\B_int[13] ), 
            .\m_cablesIn[24][13] (\m_cablesIn[24] [13]), .\B_int[14] (\B_int[14] ), 
            .\m_cablesIn[24][14] (\m_cablesIn[24] [14]), .\m_cablesIn[25][14] (\m_cablesIn[25] [14]), 
            .\m_cablesIn[25][15] (\m_cablesIn[25] [15]), .\B_int[11] (\B_int[11] ), 
            .\m_cablesIn[24][11] (\m_cablesIn[24] [11]), .\B_int[12] (\B_int[12] ), 
            .\m_cablesIn[24][12] (\m_cablesIn[24] [12]), .\m_cablesIn[25][12] (\m_cablesIn[25] [12]), 
            .\m_cablesIn[25][13] (\m_cablesIn[25] [13]), .\B_int[9] (\B_int[9] ), 
            .\m_cablesIn[24][9] (\m_cablesIn[24] [9]), .\B_int[10] (\B_int[10] ), 
            .\m_cablesIn[24][10] (\m_cablesIn[24] [10]), .\m_cablesIn[25][10] (\m_cablesIn[25] [10]), 
            .\m_cablesIn[25][11] (\m_cablesIn[25] [11]), .\B_int[7] (\B_int[7] ), 
            .\m_cablesIn[24][7] (\m_cablesIn[24] [7]), .\B_int[8] (\B_int[8] ), 
            .\m_cablesIn[24][8] (\m_cablesIn[24] [8]), .\m_cablesIn[25][8] (\m_cablesIn[25] [8]), 
            .\m_cablesIn[25][9] (\m_cablesIn[25] [9]), .\B_int[5] (\B_int[5] ), 
            .\m_cablesIn[24][5] (\m_cablesIn[24] [5]), .\B_int[6] (\B_int[6] ), 
            .\m_cablesIn[24][6] (\m_cablesIn[24] [6]), .\m_cablesIn[25][6] (\m_cablesIn[25] [6]), 
            .\m_cablesIn[25][7] (\m_cablesIn[25] [7]), .\B_int[3] (\B_int[3] ), 
            .\m_cablesIn[24][3] (\m_cablesIn[24] [3]), .\B_int[4] (\B_int[4] ), 
            .\m_cablesIn[24][4] (\m_cablesIn[24] [4]), .\m_cablesIn[25][4] (\m_cablesIn[25] [4]), 
            .\m_cablesIn[25][5] (\m_cablesIn[25] [5]), .\B_int[1] (\B_int[1] ), 
            .\m_cablesIn[24][1] (\m_cablesIn[24] [1]), .\B_int[2] (\B_int[2] ), 
            .\m_cablesIn[24][2] (\m_cablesIn[24] [2]), .\m_cablesIn[25][2] (\m_cablesIn[25] [2]), 
            .\m_cablesIn[25][3] (\m_cablesIn[25] [3]), .\B_int[0] (\B_int[0] ), 
            .\frac_div[3] (frac_div[3]), .\m_cablesIn[25][1] (\m_cablesIn[25] [1]));
    \a_s(24)_U9  \divisor_24..int_mod  (.\m_cablesIn[23][23] (\m_cablesIn[23] [23]), 
            .\QQ_in[23][22] (\QQ_in[23][22] ), .GND_net(GND_net), .\m_cablesIn[23][24] (\m_cablesIn[23] [24]), 
            .\m_cablesIn[24][24] (\m_cablesIn[24] [24]), .\QQ_in[24][23] (\QQ_in[24][23] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[23][21] (\m_cablesIn[23] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[23][22] (\m_cablesIn[23] [22]), 
            .\m_cablesIn[24][22] (\m_cablesIn[24] [22]), .\m_cablesIn[24][23] (\m_cablesIn[24] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[23][19] (\m_cablesIn[23] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[23][20] (\m_cablesIn[23] [20]), 
            .\m_cablesIn[24][20] (\m_cablesIn[24] [20]), .\m_cablesIn[24][21] (\m_cablesIn[24] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[23][17] (\m_cablesIn[23] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[23][18] (\m_cablesIn[23] [18]), 
            .\m_cablesIn[24][18] (\m_cablesIn[24] [18]), .\m_cablesIn[24][19] (\m_cablesIn[24] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[23][15] (\m_cablesIn[23] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[23][16] (\m_cablesIn[23] [16]), 
            .\m_cablesIn[24][16] (\m_cablesIn[24] [16]), .\m_cablesIn[24][17] (\m_cablesIn[24] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[23][13] (\m_cablesIn[23] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[23][14] (\m_cablesIn[23] [14]), 
            .\m_cablesIn[24][14] (\m_cablesIn[24] [14]), .\m_cablesIn[24][15] (\m_cablesIn[24] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[23][11] (\m_cablesIn[23] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[23][12] (\m_cablesIn[23] [12]), 
            .\m_cablesIn[24][12] (\m_cablesIn[24] [12]), .\m_cablesIn[24][13] (\m_cablesIn[24] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[23][9] (\m_cablesIn[23] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[23][10] (\m_cablesIn[23] [10]), 
            .\m_cablesIn[24][10] (\m_cablesIn[24] [10]), .\m_cablesIn[24][11] (\m_cablesIn[24] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[23][7] (\m_cablesIn[23] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[23][8] (\m_cablesIn[23] [8]), 
            .\m_cablesIn[24][8] (\m_cablesIn[24] [8]), .\m_cablesIn[24][9] (\m_cablesIn[24] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[23][5] (\m_cablesIn[23] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[23][6] (\m_cablesIn[23] [6]), 
            .\m_cablesIn[24][6] (\m_cablesIn[24] [6]), .\m_cablesIn[24][7] (\m_cablesIn[24] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[23][3] (\m_cablesIn[23] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[23][4] (\m_cablesIn[23] [4]), 
            .\m_cablesIn[24][4] (\m_cablesIn[24] [4]), .\m_cablesIn[24][5] (\m_cablesIn[24] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[23][1] (\m_cablesIn[23] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[23][2] (\m_cablesIn[23] [2]), 
            .\m_cablesIn[24][2] (\m_cablesIn[24] [2]), .\m_cablesIn[24][3] (\m_cablesIn[24] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[4] (frac_div[4]), .\m_cablesIn[24][1] (\m_cablesIn[24] [1]));
    \a_s(24)_U10  \divisor_23..int_mod  (.\m_cablesIn[22][23] (\m_cablesIn[22] [23]), 
            .\QQ_in[22][21] (\QQ_in[22][21] ), .GND_net(GND_net), .\m_cablesIn[22][24] (\m_cablesIn[22] [24]), 
            .\m_cablesIn[23][24] (\m_cablesIn[23] [24]), .\QQ_in[23][22] (\QQ_in[23][22] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[22][21] (\m_cablesIn[22] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[22][22] (\m_cablesIn[22] [22]), 
            .\m_cablesIn[23][22] (\m_cablesIn[23] [22]), .\m_cablesIn[23][23] (\m_cablesIn[23] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[22][19] (\m_cablesIn[22] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[22][20] (\m_cablesIn[22] [20]), 
            .\m_cablesIn[23][20] (\m_cablesIn[23] [20]), .\m_cablesIn[23][21] (\m_cablesIn[23] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[22][17] (\m_cablesIn[22] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[22][18] (\m_cablesIn[22] [18]), 
            .\m_cablesIn[23][18] (\m_cablesIn[23] [18]), .\m_cablesIn[23][19] (\m_cablesIn[23] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[22][15] (\m_cablesIn[22] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[22][16] (\m_cablesIn[22] [16]), 
            .\m_cablesIn[23][16] (\m_cablesIn[23] [16]), .\m_cablesIn[23][17] (\m_cablesIn[23] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[22][13] (\m_cablesIn[22] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[22][14] (\m_cablesIn[22] [14]), 
            .\m_cablesIn[23][14] (\m_cablesIn[23] [14]), .\m_cablesIn[23][15] (\m_cablesIn[23] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[22][11] (\m_cablesIn[22] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[22][12] (\m_cablesIn[22] [12]), 
            .\m_cablesIn[23][12] (\m_cablesIn[23] [12]), .\m_cablesIn[23][13] (\m_cablesIn[23] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[22][9] (\m_cablesIn[22] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[22][10] (\m_cablesIn[22] [10]), 
            .\m_cablesIn[23][10] (\m_cablesIn[23] [10]), .\m_cablesIn[23][11] (\m_cablesIn[23] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[22][7] (\m_cablesIn[22] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[22][8] (\m_cablesIn[22] [8]), 
            .\m_cablesIn[23][8] (\m_cablesIn[23] [8]), .\m_cablesIn[23][9] (\m_cablesIn[23] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[22][5] (\m_cablesIn[22] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[22][6] (\m_cablesIn[22] [6]), 
            .\m_cablesIn[23][6] (\m_cablesIn[23] [6]), .\m_cablesIn[23][7] (\m_cablesIn[23] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[22][3] (\m_cablesIn[22] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[22][4] (\m_cablesIn[22] [4]), 
            .\m_cablesIn[23][4] (\m_cablesIn[23] [4]), .\m_cablesIn[23][5] (\m_cablesIn[23] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[22][1] (\m_cablesIn[22] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[22][2] (\m_cablesIn[22] [2]), 
            .\m_cablesIn[23][2] (\m_cablesIn[23] [2]), .\m_cablesIn[23][3] (\m_cablesIn[23] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[5] (frac_div[5]), .\m_cablesIn[23][1] (\m_cablesIn[23] [1]));
    \a_s(24)_U11  \divisor_22..int_mod  (.\m_cablesIn[21][23] (\m_cablesIn[21] [23]), 
            .\QQ_in[21][20] (\QQ_in[21][20] ), .GND_net(GND_net), .\m_cablesIn[21][24] (\m_cablesIn[21] [24]), 
            .\m_cablesIn[22][24] (\m_cablesIn[22] [24]), .\QQ_in[22][21] (\QQ_in[22][21] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[21][21] (\m_cablesIn[21] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[21][22] (\m_cablesIn[21] [22]), 
            .\m_cablesIn[22][22] (\m_cablesIn[22] [22]), .\m_cablesIn[22][23] (\m_cablesIn[22] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[21][19] (\m_cablesIn[21] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[21][20] (\m_cablesIn[21] [20]), 
            .\m_cablesIn[22][20] (\m_cablesIn[22] [20]), .\m_cablesIn[22][21] (\m_cablesIn[22] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[21][17] (\m_cablesIn[21] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[21][18] (\m_cablesIn[21] [18]), 
            .\m_cablesIn[22][18] (\m_cablesIn[22] [18]), .\m_cablesIn[22][19] (\m_cablesIn[22] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[21][15] (\m_cablesIn[21] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[21][16] (\m_cablesIn[21] [16]), 
            .\m_cablesIn[22][16] (\m_cablesIn[22] [16]), .\m_cablesIn[22][17] (\m_cablesIn[22] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[21][13] (\m_cablesIn[21] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[21][14] (\m_cablesIn[21] [14]), 
            .\m_cablesIn[22][14] (\m_cablesIn[22] [14]), .\m_cablesIn[22][15] (\m_cablesIn[22] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[21][11] (\m_cablesIn[21] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[21][12] (\m_cablesIn[21] [12]), 
            .\m_cablesIn[22][12] (\m_cablesIn[22] [12]), .\m_cablesIn[22][13] (\m_cablesIn[22] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[21][9] (\m_cablesIn[21] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[21][10] (\m_cablesIn[21] [10]), 
            .\m_cablesIn[22][10] (\m_cablesIn[22] [10]), .\m_cablesIn[22][11] (\m_cablesIn[22] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[21][7] (\m_cablesIn[21] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[21][8] (\m_cablesIn[21] [8]), 
            .\m_cablesIn[22][8] (\m_cablesIn[22] [8]), .\m_cablesIn[22][9] (\m_cablesIn[22] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[21][5] (\m_cablesIn[21] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[21][6] (\m_cablesIn[21] [6]), 
            .\m_cablesIn[22][6] (\m_cablesIn[22] [6]), .\m_cablesIn[22][7] (\m_cablesIn[22] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[21][3] (\m_cablesIn[21] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[21][4] (\m_cablesIn[21] [4]), 
            .\m_cablesIn[22][4] (\m_cablesIn[22] [4]), .\m_cablesIn[22][5] (\m_cablesIn[22] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[21][1] (\m_cablesIn[21] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[21][2] (\m_cablesIn[21] [2]), 
            .\m_cablesIn[22][2] (\m_cablesIn[22] [2]), .\m_cablesIn[22][3] (\m_cablesIn[22] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[6] (frac_div[6]), .\m_cablesIn[22][1] (\m_cablesIn[22] [1]));
    \a_s(24)_U12  \divisor_21..int_mod  (.\m_cablesIn[20][23] (\m_cablesIn[20] [23]), 
            .\QQ_in[20][19] (\QQ_in[20][19] ), .GND_net(GND_net), .\m_cablesIn[20][24] (\m_cablesIn[20] [24]), 
            .\m_cablesIn[21][24] (\m_cablesIn[21] [24]), .\QQ_in[21][20] (\QQ_in[21][20] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[20][21] (\m_cablesIn[20] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[20][22] (\m_cablesIn[20] [22]), 
            .\m_cablesIn[21][22] (\m_cablesIn[21] [22]), .\m_cablesIn[21][23] (\m_cablesIn[21] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[20][19] (\m_cablesIn[20] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[20][20] (\m_cablesIn[20] [20]), 
            .\m_cablesIn[21][20] (\m_cablesIn[21] [20]), .\m_cablesIn[21][21] (\m_cablesIn[21] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[20][17] (\m_cablesIn[20] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[20][18] (\m_cablesIn[20] [18]), 
            .\m_cablesIn[21][18] (\m_cablesIn[21] [18]), .\m_cablesIn[21][19] (\m_cablesIn[21] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[20][15] (\m_cablesIn[20] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[20][16] (\m_cablesIn[20] [16]), 
            .\m_cablesIn[21][16] (\m_cablesIn[21] [16]), .\m_cablesIn[21][17] (\m_cablesIn[21] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[20][13] (\m_cablesIn[20] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[20][14] (\m_cablesIn[20] [14]), 
            .\m_cablesIn[21][14] (\m_cablesIn[21] [14]), .\m_cablesIn[21][15] (\m_cablesIn[21] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[20][11] (\m_cablesIn[20] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[20][12] (\m_cablesIn[20] [12]), 
            .\m_cablesIn[21][12] (\m_cablesIn[21] [12]), .\m_cablesIn[21][13] (\m_cablesIn[21] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[20][9] (\m_cablesIn[20] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[20][10] (\m_cablesIn[20] [10]), 
            .\m_cablesIn[21][10] (\m_cablesIn[21] [10]), .\m_cablesIn[21][11] (\m_cablesIn[21] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[20][7] (\m_cablesIn[20] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[20][8] (\m_cablesIn[20] [8]), 
            .\m_cablesIn[21][8] (\m_cablesIn[21] [8]), .\m_cablesIn[21][9] (\m_cablesIn[21] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[20][5] (\m_cablesIn[20] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[20][6] (\m_cablesIn[20] [6]), 
            .\m_cablesIn[21][6] (\m_cablesIn[21] [6]), .\m_cablesIn[21][7] (\m_cablesIn[21] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[20][3] (\m_cablesIn[20] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[20][4] (\m_cablesIn[20] [4]), 
            .\m_cablesIn[21][4] (\m_cablesIn[21] [4]), .\m_cablesIn[21][5] (\m_cablesIn[21] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[20][1] (\m_cablesIn[20] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[20][2] (\m_cablesIn[20] [2]), 
            .\m_cablesIn[21][2] (\m_cablesIn[21] [2]), .\m_cablesIn[21][3] (\m_cablesIn[21] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[7] (frac_div[7]), .\m_cablesIn[21][1] (\m_cablesIn[21] [1]));
    \a_s(24)_U13  \divisor_20..int_mod  (.\m_cablesIn[19][23] (\m_cablesIn[19] [23]), 
            .\QQ_in[19][18] (\QQ_in[19][18] ), .GND_net(GND_net), .\m_cablesIn[19][24] (\m_cablesIn[19] [24]), 
            .\m_cablesIn[20][24] (\m_cablesIn[20] [24]), .\QQ_in[20][19] (\QQ_in[20][19] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[19][21] (\m_cablesIn[19] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[19][22] (\m_cablesIn[19] [22]), 
            .\m_cablesIn[20][22] (\m_cablesIn[20] [22]), .\m_cablesIn[20][23] (\m_cablesIn[20] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[19][19] (\m_cablesIn[19] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[19][20] (\m_cablesIn[19] [20]), 
            .\m_cablesIn[20][20] (\m_cablesIn[20] [20]), .\m_cablesIn[20][21] (\m_cablesIn[20] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[19][17] (\m_cablesIn[19] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[19][18] (\m_cablesIn[19] [18]), 
            .\m_cablesIn[20][18] (\m_cablesIn[20] [18]), .\m_cablesIn[20][19] (\m_cablesIn[20] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[19][15] (\m_cablesIn[19] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[19][16] (\m_cablesIn[19] [16]), 
            .\m_cablesIn[20][16] (\m_cablesIn[20] [16]), .\m_cablesIn[20][17] (\m_cablesIn[20] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[19][13] (\m_cablesIn[19] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[19][14] (\m_cablesIn[19] [14]), 
            .\m_cablesIn[20][14] (\m_cablesIn[20] [14]), .\m_cablesIn[20][15] (\m_cablesIn[20] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[19][11] (\m_cablesIn[19] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[19][12] (\m_cablesIn[19] [12]), 
            .\m_cablesIn[20][12] (\m_cablesIn[20] [12]), .\m_cablesIn[20][13] (\m_cablesIn[20] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[19][9] (\m_cablesIn[19] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[19][10] (\m_cablesIn[19] [10]), 
            .\m_cablesIn[20][10] (\m_cablesIn[20] [10]), .\m_cablesIn[20][11] (\m_cablesIn[20] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[19][7] (\m_cablesIn[19] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[19][8] (\m_cablesIn[19] [8]), 
            .\m_cablesIn[20][8] (\m_cablesIn[20] [8]), .\m_cablesIn[20][9] (\m_cablesIn[20] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[19][5] (\m_cablesIn[19] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[19][6] (\m_cablesIn[19] [6]), 
            .\m_cablesIn[20][6] (\m_cablesIn[20] [6]), .\m_cablesIn[20][7] (\m_cablesIn[20] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[19][3] (\m_cablesIn[19] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[19][4] (\m_cablesIn[19] [4]), 
            .\m_cablesIn[20][4] (\m_cablesIn[20] [4]), .\m_cablesIn[20][5] (\m_cablesIn[20] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[19][1] (\m_cablesIn[19] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[19][2] (\m_cablesIn[19] [2]), 
            .\m_cablesIn[20][2] (\m_cablesIn[20] [2]), .\m_cablesIn[20][3] (\m_cablesIn[20] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[8] (frac_div[8]), .\m_cablesIn[20][1] (\m_cablesIn[20] [1]));
    \a_s(24)_U14  \divisor_1..int_mod  (.GND_net(GND_net), .\m_cablesIn[1][24] (\m_cablesIn[1] [24]), 
            .\QQ_in[1][0] (\QQ_in[1][0] ), .\A_int[21] (\A_int[21] ), .\B_int[21] (\B_int[21] ), 
            .\A_int[22] (\A_int[22] ), .\B_int[22] (\B_int[22] ), .\m_cablesIn[1][22] (\m_cablesIn[1] [22]), 
            .\m_cablesIn[1][23] (\m_cablesIn[1] [23]), .\A_int[19] (\A_int[19] ), 
            .\B_int[19] (\B_int[19] ), .\A_int[20] (\A_int[20] ), .\B_int[20] (\B_int[20] ), 
            .\m_cablesIn[1][20] (\m_cablesIn[1] [20]), .\m_cablesIn[1][21] (\m_cablesIn[1] [21]), 
            .\A_int[17] (\A_int[17] ), .\B_int[17] (\B_int[17] ), .\A_int[18] (\A_int[18] ), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[1][18] (\m_cablesIn[1] [18]), 
            .\m_cablesIn[1][19] (\m_cablesIn[1] [19]), .\A_int[15] (\A_int[15] ), 
            .\B_int[15] (\B_int[15] ), .\A_int[16] (\A_int[16] ), .\B_int[16] (\B_int[16] ), 
            .\m_cablesIn[1][16] (\m_cablesIn[1] [16]), .\m_cablesIn[1][17] (\m_cablesIn[1] [17]), 
            .\A_int[13] (\A_int[13] ), .\B_int[13] (\B_int[13] ), .\A_int[14] (\A_int[14] ), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[1][14] (\m_cablesIn[1] [14]), 
            .\m_cablesIn[1][15] (\m_cablesIn[1] [15]), .\A_int[11] (\A_int[11] ), 
            .\B_int[11] (\B_int[11] ), .\A_int[12] (\A_int[12] ), .\B_int[12] (\B_int[12] ), 
            .\m_cablesIn[1][12] (\m_cablesIn[1] [12]), .\m_cablesIn[1][13] (\m_cablesIn[1] [13]), 
            .\A_int[9] (\A_int[9] ), .\B_int[9] (\B_int[9] ), .\A_int[10] (\A_int[10] ), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[1][10] (\m_cablesIn[1] [10]), 
            .\m_cablesIn[1][11] (\m_cablesIn[1] [11]), .\A_int[7] (\A_int[7] ), 
            .\B_int[7] (\B_int[7] ), .\A_int[8] (\A_int[8] ), .\B_int[8] (\B_int[8] ), 
            .\m_cablesIn[1][8] (\m_cablesIn[1] [8]), .\m_cablesIn[1][9] (\m_cablesIn[1] [9]), 
            .\A_int[5] (\A_int[5] ), .\B_int[5] (\B_int[5] ), .\A_int[6] (\A_int[6] ), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[1][6] (\m_cablesIn[1] [6]), 
            .\m_cablesIn[1][7] (\m_cablesIn[1] [7]), .\A_int[3] (\A_int[3] ), 
            .\B_int[3] (\B_int[3] ), .\A_int[4] (\A_int[4] ), .\B_int[4] (\B_int[4] ), 
            .\m_cablesIn[1][4] (\m_cablesIn[1] [4]), .\m_cablesIn[1][5] (\m_cablesIn[1] [5]), 
            .\A_int[1] (\A_int[1] ), .\B_int[1] (\B_int[1] ), .\A_int[2] (\A_int[2] ), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[1][2] (\m_cablesIn[1] [2]), 
            .\m_cablesIn[1][3] (\m_cablesIn[1] [3]), .\A_int[0] (\A_int[0] ), 
            .\B_int[0] (\B_int[0] ), .\m_cablesIn[1][1] (\m_cablesIn[1] [1]));
    \a_s(24)_U15  \divisor_19..int_mod  (.\m_cablesIn[18][23] (\m_cablesIn[18] [23]), 
            .\QQ_in[18][17] (\QQ_in[18][17] ), .GND_net(GND_net), .\m_cablesIn[18][24] (\m_cablesIn[18] [24]), 
            .\m_cablesIn[19][24] (\m_cablesIn[19] [24]), .\QQ_in[19][18] (\QQ_in[19][18] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[18][21] (\m_cablesIn[18] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[18][22] (\m_cablesIn[18] [22]), 
            .\m_cablesIn[19][22] (\m_cablesIn[19] [22]), .\m_cablesIn[19][23] (\m_cablesIn[19] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[18][19] (\m_cablesIn[18] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[18][20] (\m_cablesIn[18] [20]), 
            .\m_cablesIn[19][20] (\m_cablesIn[19] [20]), .\m_cablesIn[19][21] (\m_cablesIn[19] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[18][17] (\m_cablesIn[18] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[18][18] (\m_cablesIn[18] [18]), 
            .\m_cablesIn[19][18] (\m_cablesIn[19] [18]), .\m_cablesIn[19][19] (\m_cablesIn[19] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[18][15] (\m_cablesIn[18] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[18][16] (\m_cablesIn[18] [16]), 
            .\m_cablesIn[19][16] (\m_cablesIn[19] [16]), .\m_cablesIn[19][17] (\m_cablesIn[19] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[18][13] (\m_cablesIn[18] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[18][14] (\m_cablesIn[18] [14]), 
            .\m_cablesIn[19][14] (\m_cablesIn[19] [14]), .\m_cablesIn[19][15] (\m_cablesIn[19] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[18][11] (\m_cablesIn[18] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[18][12] (\m_cablesIn[18] [12]), 
            .\m_cablesIn[19][12] (\m_cablesIn[19] [12]), .\m_cablesIn[19][13] (\m_cablesIn[19] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[18][9] (\m_cablesIn[18] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[18][10] (\m_cablesIn[18] [10]), 
            .\m_cablesIn[19][10] (\m_cablesIn[19] [10]), .\m_cablesIn[19][11] (\m_cablesIn[19] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[18][7] (\m_cablesIn[18] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[18][8] (\m_cablesIn[18] [8]), 
            .\m_cablesIn[19][8] (\m_cablesIn[19] [8]), .\m_cablesIn[19][9] (\m_cablesIn[19] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[18][5] (\m_cablesIn[18] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[18][6] (\m_cablesIn[18] [6]), 
            .\m_cablesIn[19][6] (\m_cablesIn[19] [6]), .\m_cablesIn[19][7] (\m_cablesIn[19] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[18][3] (\m_cablesIn[18] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[18][4] (\m_cablesIn[18] [4]), 
            .\m_cablesIn[19][4] (\m_cablesIn[19] [4]), .\m_cablesIn[19][5] (\m_cablesIn[19] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[18][1] (\m_cablesIn[18] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[18][2] (\m_cablesIn[18] [2]), 
            .\m_cablesIn[19][2] (\m_cablesIn[19] [2]), .\m_cablesIn[19][3] (\m_cablesIn[19] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[9] (frac_div[9]), .\m_cablesIn[19][1] (\m_cablesIn[19] [1]));
    \a_s(24)_U16  \divisor_18..int_mod  (.\m_cablesIn[17][23] (\m_cablesIn[17] [23]), 
            .\QQ_in[17][16] (\QQ_in[17][16] ), .GND_net(GND_net), .\m_cablesIn[17][24] (\m_cablesIn[17] [24]), 
            .\m_cablesIn[18][24] (\m_cablesIn[18] [24]), .\QQ_in[18][17] (\QQ_in[18][17] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[17][21] (\m_cablesIn[17] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[17][22] (\m_cablesIn[17] [22]), 
            .\m_cablesIn[18][22] (\m_cablesIn[18] [22]), .\m_cablesIn[18][23] (\m_cablesIn[18] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[17][19] (\m_cablesIn[17] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[17][20] (\m_cablesIn[17] [20]), 
            .\m_cablesIn[18][20] (\m_cablesIn[18] [20]), .\m_cablesIn[18][21] (\m_cablesIn[18] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[17][17] (\m_cablesIn[17] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[17][18] (\m_cablesIn[17] [18]), 
            .\m_cablesIn[18][18] (\m_cablesIn[18] [18]), .\m_cablesIn[18][19] (\m_cablesIn[18] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[17][15] (\m_cablesIn[17] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[17][16] (\m_cablesIn[17] [16]), 
            .\m_cablesIn[18][16] (\m_cablesIn[18] [16]), .\m_cablesIn[18][17] (\m_cablesIn[18] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[17][13] (\m_cablesIn[17] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[17][14] (\m_cablesIn[17] [14]), 
            .\m_cablesIn[18][14] (\m_cablesIn[18] [14]), .\m_cablesIn[18][15] (\m_cablesIn[18] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[17][11] (\m_cablesIn[17] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[17][12] (\m_cablesIn[17] [12]), 
            .\m_cablesIn[18][12] (\m_cablesIn[18] [12]), .\m_cablesIn[18][13] (\m_cablesIn[18] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[17][9] (\m_cablesIn[17] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[17][10] (\m_cablesIn[17] [10]), 
            .\m_cablesIn[18][10] (\m_cablesIn[18] [10]), .\m_cablesIn[18][11] (\m_cablesIn[18] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[17][7] (\m_cablesIn[17] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[17][8] (\m_cablesIn[17] [8]), 
            .\m_cablesIn[18][8] (\m_cablesIn[18] [8]), .\m_cablesIn[18][9] (\m_cablesIn[18] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[17][5] (\m_cablesIn[17] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[17][6] (\m_cablesIn[17] [6]), 
            .\m_cablesIn[18][6] (\m_cablesIn[18] [6]), .\m_cablesIn[18][7] (\m_cablesIn[18] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[17][3] (\m_cablesIn[17] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[17][4] (\m_cablesIn[17] [4]), 
            .\m_cablesIn[18][4] (\m_cablesIn[18] [4]), .\m_cablesIn[18][5] (\m_cablesIn[18] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[17][1] (\m_cablesIn[17] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[17][2] (\m_cablesIn[17] [2]), 
            .\m_cablesIn[18][2] (\m_cablesIn[18] [2]), .\m_cablesIn[18][3] (\m_cablesIn[18] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[10] (frac_div[10]), .\m_cablesIn[18][1] (\m_cablesIn[18] [1]));
    \a_s(24)_U17  \divisor_17..int_mod  (.\m_cablesIn[16][23] (\m_cablesIn[16] [23]), 
            .\QQ_in[16][15] (\QQ_in[16][15] ), .GND_net(GND_net), .\m_cablesIn[16][24] (\m_cablesIn[16] [24]), 
            .\m_cablesIn[17][24] (\m_cablesIn[17] [24]), .\QQ_in[17][16] (\QQ_in[17][16] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[16][21] (\m_cablesIn[16] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[16][22] (\m_cablesIn[16] [22]), 
            .\m_cablesIn[17][22] (\m_cablesIn[17] [22]), .\m_cablesIn[17][23] (\m_cablesIn[17] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[16][19] (\m_cablesIn[16] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[16][20] (\m_cablesIn[16] [20]), 
            .\m_cablesIn[17][20] (\m_cablesIn[17] [20]), .\m_cablesIn[17][21] (\m_cablesIn[17] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[16][17] (\m_cablesIn[16] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[16][18] (\m_cablesIn[16] [18]), 
            .\m_cablesIn[17][18] (\m_cablesIn[17] [18]), .\m_cablesIn[17][19] (\m_cablesIn[17] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[16][15] (\m_cablesIn[16] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[16][16] (\m_cablesIn[16] [16]), 
            .\m_cablesIn[17][16] (\m_cablesIn[17] [16]), .\m_cablesIn[17][17] (\m_cablesIn[17] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[16][13] (\m_cablesIn[16] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[16][14] (\m_cablesIn[16] [14]), 
            .\m_cablesIn[17][14] (\m_cablesIn[17] [14]), .\m_cablesIn[17][15] (\m_cablesIn[17] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[16][11] (\m_cablesIn[16] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[16][12] (\m_cablesIn[16] [12]), 
            .\m_cablesIn[17][12] (\m_cablesIn[17] [12]), .\m_cablesIn[17][13] (\m_cablesIn[17] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[16][9] (\m_cablesIn[16] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[16][10] (\m_cablesIn[16] [10]), 
            .\m_cablesIn[17][10] (\m_cablesIn[17] [10]), .\m_cablesIn[17][11] (\m_cablesIn[17] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[16][7] (\m_cablesIn[16] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[16][8] (\m_cablesIn[16] [8]), 
            .\m_cablesIn[17][8] (\m_cablesIn[17] [8]), .\m_cablesIn[17][9] (\m_cablesIn[17] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[16][5] (\m_cablesIn[16] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[16][6] (\m_cablesIn[16] [6]), 
            .\m_cablesIn[17][6] (\m_cablesIn[17] [6]), .\m_cablesIn[17][7] (\m_cablesIn[17] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[16][3] (\m_cablesIn[16] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[16][4] (\m_cablesIn[16] [4]), 
            .\m_cablesIn[17][4] (\m_cablesIn[17] [4]), .\m_cablesIn[17][5] (\m_cablesIn[17] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[16][1] (\m_cablesIn[16] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[16][2] (\m_cablesIn[16] [2]), 
            .\m_cablesIn[17][2] (\m_cablesIn[17] [2]), .\m_cablesIn[17][3] (\m_cablesIn[17] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[11] (frac_div[11]), .\m_cablesIn[17][1] (\m_cablesIn[17] [1]));
    \a_s(24)_U18  \divisor_16..int_mod  (.\m_cablesIn[15][23] (\m_cablesIn[15] [23]), 
            .\QQ_in[15][14] (\QQ_in[15][14] ), .GND_net(GND_net), .\m_cablesIn[15][24] (\m_cablesIn[15] [24]), 
            .\m_cablesIn[16][24] (\m_cablesIn[16] [24]), .\QQ_in[16][15] (\QQ_in[16][15] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[15][21] (\m_cablesIn[15] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[15][22] (\m_cablesIn[15] [22]), 
            .\m_cablesIn[16][22] (\m_cablesIn[16] [22]), .\m_cablesIn[16][23] (\m_cablesIn[16] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[15][19] (\m_cablesIn[15] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[15][20] (\m_cablesIn[15] [20]), 
            .\m_cablesIn[16][20] (\m_cablesIn[16] [20]), .\m_cablesIn[16][21] (\m_cablesIn[16] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[15][17] (\m_cablesIn[15] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[15][18] (\m_cablesIn[15] [18]), 
            .\m_cablesIn[16][18] (\m_cablesIn[16] [18]), .\m_cablesIn[16][19] (\m_cablesIn[16] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[15][15] (\m_cablesIn[15] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[15][16] (\m_cablesIn[15] [16]), 
            .\m_cablesIn[16][16] (\m_cablesIn[16] [16]), .\m_cablesIn[16][17] (\m_cablesIn[16] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[15][13] (\m_cablesIn[15] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[15][14] (\m_cablesIn[15] [14]), 
            .\m_cablesIn[16][14] (\m_cablesIn[16] [14]), .\m_cablesIn[16][15] (\m_cablesIn[16] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[15][11] (\m_cablesIn[15] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[15][12] (\m_cablesIn[15] [12]), 
            .\m_cablesIn[16][12] (\m_cablesIn[16] [12]), .\m_cablesIn[16][13] (\m_cablesIn[16] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[15][9] (\m_cablesIn[15] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[15][10] (\m_cablesIn[15] [10]), 
            .\m_cablesIn[16][10] (\m_cablesIn[16] [10]), .\m_cablesIn[16][11] (\m_cablesIn[16] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[15][7] (\m_cablesIn[15] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[15][8] (\m_cablesIn[15] [8]), 
            .\m_cablesIn[16][8] (\m_cablesIn[16] [8]), .\m_cablesIn[16][9] (\m_cablesIn[16] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[15][5] (\m_cablesIn[15] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[15][6] (\m_cablesIn[15] [6]), 
            .\m_cablesIn[16][6] (\m_cablesIn[16] [6]), .\m_cablesIn[16][7] (\m_cablesIn[16] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[15][3] (\m_cablesIn[15] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[15][4] (\m_cablesIn[15] [4]), 
            .\m_cablesIn[16][4] (\m_cablesIn[16] [4]), .\m_cablesIn[16][5] (\m_cablesIn[16] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[15][1] (\m_cablesIn[15] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[15][2] (\m_cablesIn[15] [2]), 
            .\m_cablesIn[16][2] (\m_cablesIn[16] [2]), .\m_cablesIn[16][3] (\m_cablesIn[16] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[12] (frac_div[12]), .\m_cablesIn[16][1] (\m_cablesIn[16] [1]));
    \a_s(24)_U19  \divisor_15..int_mod  (.\m_cablesIn[14][23] (\m_cablesIn[14] [23]), 
            .\QQ_in[14][13] (\QQ_in[14][13] ), .GND_net(GND_net), .\m_cablesIn[14][24] (\m_cablesIn[14] [24]), 
            .\m_cablesIn[15][24] (\m_cablesIn[15] [24]), .\QQ_in[15][14] (\QQ_in[15][14] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[14][21] (\m_cablesIn[14] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[14][22] (\m_cablesIn[14] [22]), 
            .\m_cablesIn[15][22] (\m_cablesIn[15] [22]), .\m_cablesIn[15][23] (\m_cablesIn[15] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[14][19] (\m_cablesIn[14] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[14][20] (\m_cablesIn[14] [20]), 
            .\m_cablesIn[15][20] (\m_cablesIn[15] [20]), .\m_cablesIn[15][21] (\m_cablesIn[15] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[14][17] (\m_cablesIn[14] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[14][18] (\m_cablesIn[14] [18]), 
            .\m_cablesIn[15][18] (\m_cablesIn[15] [18]), .\m_cablesIn[15][19] (\m_cablesIn[15] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[14][15] (\m_cablesIn[14] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[14][16] (\m_cablesIn[14] [16]), 
            .\m_cablesIn[15][16] (\m_cablesIn[15] [16]), .\m_cablesIn[15][17] (\m_cablesIn[15] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[14][13] (\m_cablesIn[14] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[14][14] (\m_cablesIn[14] [14]), 
            .\m_cablesIn[15][14] (\m_cablesIn[15] [14]), .\m_cablesIn[15][15] (\m_cablesIn[15] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[14][11] (\m_cablesIn[14] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[14][12] (\m_cablesIn[14] [12]), 
            .\m_cablesIn[15][12] (\m_cablesIn[15] [12]), .\m_cablesIn[15][13] (\m_cablesIn[15] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[14][9] (\m_cablesIn[14] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[14][10] (\m_cablesIn[14] [10]), 
            .\m_cablesIn[15][10] (\m_cablesIn[15] [10]), .\m_cablesIn[15][11] (\m_cablesIn[15] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[14][7] (\m_cablesIn[14] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[14][8] (\m_cablesIn[14] [8]), 
            .\m_cablesIn[15][8] (\m_cablesIn[15] [8]), .\m_cablesIn[15][9] (\m_cablesIn[15] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[14][5] (\m_cablesIn[14] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[14][6] (\m_cablesIn[14] [6]), 
            .\m_cablesIn[15][6] (\m_cablesIn[15] [6]), .\m_cablesIn[15][7] (\m_cablesIn[15] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[14][3] (\m_cablesIn[14] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[14][4] (\m_cablesIn[14] [4]), 
            .\m_cablesIn[15][4] (\m_cablesIn[15] [4]), .\m_cablesIn[15][5] (\m_cablesIn[15] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[14][1] (\m_cablesIn[14] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[14][2] (\m_cablesIn[14] [2]), 
            .\m_cablesIn[15][2] (\m_cablesIn[15] [2]), .\m_cablesIn[15][3] (\m_cablesIn[15] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[13] (frac_div[13]), .\m_cablesIn[15][1] (\m_cablesIn[15] [1]));
    \a_s(24)_U20  \divisor_14..int_mod  (.\m_cablesIn[13][23] (\m_cablesIn[13] [23]), 
            .\QQ_in[13][12] (\QQ_in[13][12] ), .GND_net(GND_net), .\m_cablesIn[13][24] (\m_cablesIn[13] [24]), 
            .\m_cablesIn[14][24] (\m_cablesIn[14] [24]), .\QQ_in[14][13] (\QQ_in[14][13] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[13][21] (\m_cablesIn[13] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[13][22] (\m_cablesIn[13] [22]), 
            .\m_cablesIn[14][22] (\m_cablesIn[14] [22]), .\m_cablesIn[14][23] (\m_cablesIn[14] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[13][19] (\m_cablesIn[13] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[13][20] (\m_cablesIn[13] [20]), 
            .\m_cablesIn[14][20] (\m_cablesIn[14] [20]), .\m_cablesIn[14][21] (\m_cablesIn[14] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[13][17] (\m_cablesIn[13] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[13][18] (\m_cablesIn[13] [18]), 
            .\m_cablesIn[14][18] (\m_cablesIn[14] [18]), .\m_cablesIn[14][19] (\m_cablesIn[14] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[13][15] (\m_cablesIn[13] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[13][16] (\m_cablesIn[13] [16]), 
            .\m_cablesIn[14][16] (\m_cablesIn[14] [16]), .\m_cablesIn[14][17] (\m_cablesIn[14] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[13][13] (\m_cablesIn[13] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[13][14] (\m_cablesIn[13] [14]), 
            .\m_cablesIn[14][14] (\m_cablesIn[14] [14]), .\m_cablesIn[14][15] (\m_cablesIn[14] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[13][11] (\m_cablesIn[13] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[13][12] (\m_cablesIn[13] [12]), 
            .\m_cablesIn[14][12] (\m_cablesIn[14] [12]), .\m_cablesIn[14][13] (\m_cablesIn[14] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[13][9] (\m_cablesIn[13] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[13][10] (\m_cablesIn[13] [10]), 
            .\m_cablesIn[14][10] (\m_cablesIn[14] [10]), .\m_cablesIn[14][11] (\m_cablesIn[14] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[13][7] (\m_cablesIn[13] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[13][8] (\m_cablesIn[13] [8]), 
            .\m_cablesIn[14][8] (\m_cablesIn[14] [8]), .\m_cablesIn[14][9] (\m_cablesIn[14] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[13][5] (\m_cablesIn[13] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[13][6] (\m_cablesIn[13] [6]), 
            .\m_cablesIn[14][6] (\m_cablesIn[14] [6]), .\m_cablesIn[14][7] (\m_cablesIn[14] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[13][3] (\m_cablesIn[13] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[13][4] (\m_cablesIn[13] [4]), 
            .\m_cablesIn[14][4] (\m_cablesIn[14] [4]), .\m_cablesIn[14][5] (\m_cablesIn[14] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[13][1] (\m_cablesIn[13] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[13][2] (\m_cablesIn[13] [2]), 
            .\m_cablesIn[14][2] (\m_cablesIn[14] [2]), .\m_cablesIn[14][3] (\m_cablesIn[14] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[14] (frac_div[14]), .\m_cablesIn[14][1] (\m_cablesIn[14] [1]));
    \a_s(24)_U21  \divisor_13..int_mod  (.\m_cablesIn[12][23] (\m_cablesIn[12] [23]), 
            .\QQ_in[12][11] (\QQ_in[12][11] ), .GND_net(GND_net), .\m_cablesIn[12][24] (\m_cablesIn[12] [24]), 
            .\m_cablesIn[13][24] (\m_cablesIn[13] [24]), .\QQ_in[13][12] (\QQ_in[13][12] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[12][21] (\m_cablesIn[12] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[12][22] (\m_cablesIn[12] [22]), 
            .\m_cablesIn[13][22] (\m_cablesIn[13] [22]), .\m_cablesIn[13][23] (\m_cablesIn[13] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[12][19] (\m_cablesIn[12] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[12][20] (\m_cablesIn[12] [20]), 
            .\m_cablesIn[13][20] (\m_cablesIn[13] [20]), .\m_cablesIn[13][21] (\m_cablesIn[13] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[12][17] (\m_cablesIn[12] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[12][18] (\m_cablesIn[12] [18]), 
            .\m_cablesIn[13][18] (\m_cablesIn[13] [18]), .\m_cablesIn[13][19] (\m_cablesIn[13] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[12][15] (\m_cablesIn[12] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[12][16] (\m_cablesIn[12] [16]), 
            .\m_cablesIn[13][16] (\m_cablesIn[13] [16]), .\m_cablesIn[13][17] (\m_cablesIn[13] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[12][13] (\m_cablesIn[12] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[12][14] (\m_cablesIn[12] [14]), 
            .\m_cablesIn[13][14] (\m_cablesIn[13] [14]), .\m_cablesIn[13][15] (\m_cablesIn[13] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[12][11] (\m_cablesIn[12] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[12][12] (\m_cablesIn[12] [12]), 
            .\m_cablesIn[13][12] (\m_cablesIn[13] [12]), .\m_cablesIn[13][13] (\m_cablesIn[13] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[12][9] (\m_cablesIn[12] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[12][10] (\m_cablesIn[12] [10]), 
            .\m_cablesIn[13][10] (\m_cablesIn[13] [10]), .\m_cablesIn[13][11] (\m_cablesIn[13] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[12][7] (\m_cablesIn[12] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[12][8] (\m_cablesIn[12] [8]), 
            .\m_cablesIn[13][8] (\m_cablesIn[13] [8]), .\m_cablesIn[13][9] (\m_cablesIn[13] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[12][5] (\m_cablesIn[12] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[12][6] (\m_cablesIn[12] [6]), 
            .\m_cablesIn[13][6] (\m_cablesIn[13] [6]), .\m_cablesIn[13][7] (\m_cablesIn[13] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[12][3] (\m_cablesIn[12] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[12][4] (\m_cablesIn[12] [4]), 
            .\m_cablesIn[13][4] (\m_cablesIn[13] [4]), .\m_cablesIn[13][5] (\m_cablesIn[13] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[12][1] (\m_cablesIn[12] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[12][2] (\m_cablesIn[12] [2]), 
            .\m_cablesIn[13][2] (\m_cablesIn[13] [2]), .\m_cablesIn[13][3] (\m_cablesIn[13] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[15] (frac_div[15]), .\m_cablesIn[13][1] (\m_cablesIn[13] [1]));
    \a_s(24)_U22  \divisor_12..int_mod  (.\m_cablesIn[11][23] (\m_cablesIn[11] [23]), 
            .\QQ_in[11][10] (\QQ_in[11][10] ), .GND_net(GND_net), .\m_cablesIn[11][24] (\m_cablesIn[11] [24]), 
            .\m_cablesIn[12][24] (\m_cablesIn[12] [24]), .\QQ_in[12][11] (\QQ_in[12][11] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[11][21] (\m_cablesIn[11] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[11][22] (\m_cablesIn[11] [22]), 
            .\m_cablesIn[12][22] (\m_cablesIn[12] [22]), .\m_cablesIn[12][23] (\m_cablesIn[12] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[11][19] (\m_cablesIn[11] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[11][20] (\m_cablesIn[11] [20]), 
            .\m_cablesIn[12][20] (\m_cablesIn[12] [20]), .\m_cablesIn[12][21] (\m_cablesIn[12] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[11][17] (\m_cablesIn[11] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[11][18] (\m_cablesIn[11] [18]), 
            .\m_cablesIn[12][18] (\m_cablesIn[12] [18]), .\m_cablesIn[12][19] (\m_cablesIn[12] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[11][15] (\m_cablesIn[11] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[11][16] (\m_cablesIn[11] [16]), 
            .\m_cablesIn[12][16] (\m_cablesIn[12] [16]), .\m_cablesIn[12][17] (\m_cablesIn[12] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[11][13] (\m_cablesIn[11] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[11][14] (\m_cablesIn[11] [14]), 
            .\m_cablesIn[12][14] (\m_cablesIn[12] [14]), .\m_cablesIn[12][15] (\m_cablesIn[12] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[11][11] (\m_cablesIn[11] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[11][12] (\m_cablesIn[11] [12]), 
            .\m_cablesIn[12][12] (\m_cablesIn[12] [12]), .\m_cablesIn[12][13] (\m_cablesIn[12] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[11][9] (\m_cablesIn[11] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[11][10] (\m_cablesIn[11] [10]), 
            .\m_cablesIn[12][10] (\m_cablesIn[12] [10]), .\m_cablesIn[12][11] (\m_cablesIn[12] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[11][7] (\m_cablesIn[11] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[11][8] (\m_cablesIn[11] [8]), 
            .\m_cablesIn[12][8] (\m_cablesIn[12] [8]), .\m_cablesIn[12][9] (\m_cablesIn[12] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[11][5] (\m_cablesIn[11] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[11][6] (\m_cablesIn[11] [6]), 
            .\m_cablesIn[12][6] (\m_cablesIn[12] [6]), .\m_cablesIn[12][7] (\m_cablesIn[12] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[11][3] (\m_cablesIn[11] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[11][4] (\m_cablesIn[11] [4]), 
            .\m_cablesIn[12][4] (\m_cablesIn[12] [4]), .\m_cablesIn[12][5] (\m_cablesIn[12] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[11][1] (\m_cablesIn[11] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[11][2] (\m_cablesIn[11] [2]), 
            .\m_cablesIn[12][2] (\m_cablesIn[12] [2]), .\m_cablesIn[12][3] (\m_cablesIn[12] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[16] (frac_div[16]), .\m_cablesIn[12][1] (\m_cablesIn[12] [1]));
    \a_s(24)_U23  \divisor_11..int_mod  (.\m_cablesIn[10][23] (\m_cablesIn[10] [23]), 
            .\QQ_in[10][9] (\QQ_in[10][9] ), .GND_net(GND_net), .\m_cablesIn[10][24] (\m_cablesIn[10] [24]), 
            .\m_cablesIn[11][24] (\m_cablesIn[11] [24]), .\QQ_in[11][10] (\QQ_in[11][10] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[10][21] (\m_cablesIn[10] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[10][22] (\m_cablesIn[10] [22]), 
            .\m_cablesIn[11][22] (\m_cablesIn[11] [22]), .\m_cablesIn[11][23] (\m_cablesIn[11] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[10][19] (\m_cablesIn[10] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[10][20] (\m_cablesIn[10] [20]), 
            .\m_cablesIn[11][20] (\m_cablesIn[11] [20]), .\m_cablesIn[11][21] (\m_cablesIn[11] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[10][17] (\m_cablesIn[10] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[10][18] (\m_cablesIn[10] [18]), 
            .\m_cablesIn[11][18] (\m_cablesIn[11] [18]), .\m_cablesIn[11][19] (\m_cablesIn[11] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[10][15] (\m_cablesIn[10] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[10][16] (\m_cablesIn[10] [16]), 
            .\m_cablesIn[11][16] (\m_cablesIn[11] [16]), .\m_cablesIn[11][17] (\m_cablesIn[11] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[10][13] (\m_cablesIn[10] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[10][14] (\m_cablesIn[10] [14]), 
            .\m_cablesIn[11][14] (\m_cablesIn[11] [14]), .\m_cablesIn[11][15] (\m_cablesIn[11] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[10][11] (\m_cablesIn[10] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[10][12] (\m_cablesIn[10] [12]), 
            .\m_cablesIn[11][12] (\m_cablesIn[11] [12]), .\m_cablesIn[11][13] (\m_cablesIn[11] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[10][9] (\m_cablesIn[10] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[10][10] (\m_cablesIn[10] [10]), 
            .\m_cablesIn[11][10] (\m_cablesIn[11] [10]), .\m_cablesIn[11][11] (\m_cablesIn[11] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[10][7] (\m_cablesIn[10] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[10][8] (\m_cablesIn[10] [8]), 
            .\m_cablesIn[11][8] (\m_cablesIn[11] [8]), .\m_cablesIn[11][9] (\m_cablesIn[11] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[10][5] (\m_cablesIn[10] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[10][6] (\m_cablesIn[10] [6]), 
            .\m_cablesIn[11][6] (\m_cablesIn[11] [6]), .\m_cablesIn[11][7] (\m_cablesIn[11] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[10][3] (\m_cablesIn[10] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[10][4] (\m_cablesIn[10] [4]), 
            .\m_cablesIn[11][4] (\m_cablesIn[11] [4]), .\m_cablesIn[11][5] (\m_cablesIn[11] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[10][1] (\m_cablesIn[10] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[10][2] (\m_cablesIn[10] [2]), 
            .\m_cablesIn[11][2] (\m_cablesIn[11] [2]), .\m_cablesIn[11][3] (\m_cablesIn[11] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[17] (frac_div[17]), .\m_cablesIn[11][1] (\m_cablesIn[11] [1]));
    \a_s(24)_U24  \divisor_10..int_mod  (.\m_cablesIn[9][23] (\m_cablesIn[9] [23]), 
            .\QQ_in[9][8] (\QQ_in[9][8] ), .GND_net(GND_net), .\m_cablesIn[9][24] (\m_cablesIn[9] [24]), 
            .\m_cablesIn[10][24] (\m_cablesIn[10] [24]), .\QQ_in[10][9] (\QQ_in[10][9] ), 
            .\B_int[21] (\B_int[21] ), .\m_cablesIn[9][21] (\m_cablesIn[9] [21]), 
            .\B_int[22] (\B_int[22] ), .\m_cablesIn[9][22] (\m_cablesIn[9] [22]), 
            .\m_cablesIn[10][22] (\m_cablesIn[10] [22]), .\m_cablesIn[10][23] (\m_cablesIn[10] [23]), 
            .\B_int[19] (\B_int[19] ), .\m_cablesIn[9][19] (\m_cablesIn[9] [19]), 
            .\B_int[20] (\B_int[20] ), .\m_cablesIn[9][20] (\m_cablesIn[9] [20]), 
            .\m_cablesIn[10][20] (\m_cablesIn[10] [20]), .\m_cablesIn[10][21] (\m_cablesIn[10] [21]), 
            .\B_int[17] (\B_int[17] ), .\m_cablesIn[9][17] (\m_cablesIn[9] [17]), 
            .\B_int[18] (\B_int[18] ), .\m_cablesIn[9][18] (\m_cablesIn[9] [18]), 
            .\m_cablesIn[10][18] (\m_cablesIn[10] [18]), .\m_cablesIn[10][19] (\m_cablesIn[10] [19]), 
            .\B_int[15] (\B_int[15] ), .\m_cablesIn[9][15] (\m_cablesIn[9] [15]), 
            .\B_int[16] (\B_int[16] ), .\m_cablesIn[9][16] (\m_cablesIn[9] [16]), 
            .\m_cablesIn[10][16] (\m_cablesIn[10] [16]), .\m_cablesIn[10][17] (\m_cablesIn[10] [17]), 
            .\B_int[13] (\B_int[13] ), .\m_cablesIn[9][13] (\m_cablesIn[9] [13]), 
            .\B_int[14] (\B_int[14] ), .\m_cablesIn[9][14] (\m_cablesIn[9] [14]), 
            .\m_cablesIn[10][14] (\m_cablesIn[10] [14]), .\m_cablesIn[10][15] (\m_cablesIn[10] [15]), 
            .\B_int[11] (\B_int[11] ), .\m_cablesIn[9][11] (\m_cablesIn[9] [11]), 
            .\B_int[12] (\B_int[12] ), .\m_cablesIn[9][12] (\m_cablesIn[9] [12]), 
            .\m_cablesIn[10][12] (\m_cablesIn[10] [12]), .\m_cablesIn[10][13] (\m_cablesIn[10] [13]), 
            .\B_int[9] (\B_int[9] ), .\m_cablesIn[9][9] (\m_cablesIn[9] [9]), 
            .\B_int[10] (\B_int[10] ), .\m_cablesIn[9][10] (\m_cablesIn[9] [10]), 
            .\m_cablesIn[10][10] (\m_cablesIn[10] [10]), .\m_cablesIn[10][11] (\m_cablesIn[10] [11]), 
            .\B_int[7] (\B_int[7] ), .\m_cablesIn[9][7] (\m_cablesIn[9] [7]), 
            .\B_int[8] (\B_int[8] ), .\m_cablesIn[9][8] (\m_cablesIn[9] [8]), 
            .\m_cablesIn[10][8] (\m_cablesIn[10] [8]), .\m_cablesIn[10][9] (\m_cablesIn[10] [9]), 
            .\B_int[5] (\B_int[5] ), .\m_cablesIn[9][5] (\m_cablesIn[9] [5]), 
            .\B_int[6] (\B_int[6] ), .\m_cablesIn[9][6] (\m_cablesIn[9] [6]), 
            .\m_cablesIn[10][6] (\m_cablesIn[10] [6]), .\m_cablesIn[10][7] (\m_cablesIn[10] [7]), 
            .\B_int[3] (\B_int[3] ), .\m_cablesIn[9][3] (\m_cablesIn[9] [3]), 
            .\B_int[4] (\B_int[4] ), .\m_cablesIn[9][4] (\m_cablesIn[9] [4]), 
            .\m_cablesIn[10][4] (\m_cablesIn[10] [4]), .\m_cablesIn[10][5] (\m_cablesIn[10] [5]), 
            .\B_int[1] (\B_int[1] ), .\m_cablesIn[9][1] (\m_cablesIn[9] [1]), 
            .\B_int[2] (\B_int[2] ), .\m_cablesIn[9][2] (\m_cablesIn[9] [2]), 
            .\m_cablesIn[10][2] (\m_cablesIn[10] [2]), .\m_cablesIn[10][3] (\m_cablesIn[10] [3]), 
            .\B_int[0] (\B_int[0] ), .\frac_div[18] (frac_div[18]), .\m_cablesIn[10][1] (\m_cablesIn[10] [1]));
    
endmodule
//
// Verilog Description of module \a_s(24) 
//

module \a_s(24)  (\m_cablesIn[8][23] , \QQ_in[8][7] , GND_net, \m_cablesIn[8][24] , 
            \m_cablesIn[9][24] , \QQ_in[9][8] , \B_int[21] , \m_cablesIn[8][21] , 
            \B_int[22] , \m_cablesIn[8][22] , \m_cablesIn[9][22] , \m_cablesIn[9][23] , 
            \B_int[19] , \m_cablesIn[8][19] , \B_int[20] , \m_cablesIn[8][20] , 
            \m_cablesIn[9][20] , \m_cablesIn[9][21] , \B_int[17] , \m_cablesIn[8][17] , 
            \B_int[18] , \m_cablesIn[8][18] , \m_cablesIn[9][18] , \m_cablesIn[9][19] , 
            \B_int[15] , \m_cablesIn[8][15] , \B_int[16] , \m_cablesIn[8][16] , 
            \m_cablesIn[9][16] , \m_cablesIn[9][17] , \B_int[13] , \m_cablesIn[8][13] , 
            \B_int[14] , \m_cablesIn[8][14] , \m_cablesIn[9][14] , \m_cablesIn[9][15] , 
            \B_int[11] , \m_cablesIn[8][11] , \B_int[12] , \m_cablesIn[8][12] , 
            \m_cablesIn[9][12] , \m_cablesIn[9][13] , \B_int[9] , \m_cablesIn[8][9] , 
            \B_int[10] , \m_cablesIn[8][10] , \m_cablesIn[9][10] , \m_cablesIn[9][11] , 
            \B_int[7] , \m_cablesIn[8][7] , \B_int[8] , \m_cablesIn[8][8] , 
            \m_cablesIn[9][8] , \m_cablesIn[9][9] , \B_int[5] , \m_cablesIn[8][5] , 
            \B_int[6] , \m_cablesIn[8][6] , \m_cablesIn[9][6] , \m_cablesIn[9][7] , 
            \B_int[3] , \m_cablesIn[8][3] , \B_int[4] , \m_cablesIn[8][4] , 
            \m_cablesIn[9][4] , \m_cablesIn[9][5] , \B_int[1] , \m_cablesIn[8][1] , 
            \B_int[2] , \m_cablesIn[8][2] , \m_cablesIn[9][2] , \m_cablesIn[9][3] , 
            \B_int[0] , \frac_div[19] , \m_cablesIn[9][1] );
    input \m_cablesIn[8][23] ;
    input \QQ_in[8][7] ;
    input GND_net;
    input \m_cablesIn[8][24] ;
    output \m_cablesIn[9][24] ;
    output \QQ_in[9][8] ;
    input \B_int[21] ;
    input \m_cablesIn[8][21] ;
    input \B_int[22] ;
    input \m_cablesIn[8][22] ;
    output \m_cablesIn[9][22] ;
    output \m_cablesIn[9][23] ;
    input \B_int[19] ;
    input \m_cablesIn[8][19] ;
    input \B_int[20] ;
    input \m_cablesIn[8][20] ;
    output \m_cablesIn[9][20] ;
    output \m_cablesIn[9][21] ;
    input \B_int[17] ;
    input \m_cablesIn[8][17] ;
    input \B_int[18] ;
    input \m_cablesIn[8][18] ;
    output \m_cablesIn[9][18] ;
    output \m_cablesIn[9][19] ;
    input \B_int[15] ;
    input \m_cablesIn[8][15] ;
    input \B_int[16] ;
    input \m_cablesIn[8][16] ;
    output \m_cablesIn[9][16] ;
    output \m_cablesIn[9][17] ;
    input \B_int[13] ;
    input \m_cablesIn[8][13] ;
    input \B_int[14] ;
    input \m_cablesIn[8][14] ;
    output \m_cablesIn[9][14] ;
    output \m_cablesIn[9][15] ;
    input \B_int[11] ;
    input \m_cablesIn[8][11] ;
    input \B_int[12] ;
    input \m_cablesIn[8][12] ;
    output \m_cablesIn[9][12] ;
    output \m_cablesIn[9][13] ;
    input \B_int[9] ;
    input \m_cablesIn[8][9] ;
    input \B_int[10] ;
    input \m_cablesIn[8][10] ;
    output \m_cablesIn[9][10] ;
    output \m_cablesIn[9][11] ;
    input \B_int[7] ;
    input \m_cablesIn[8][7] ;
    input \B_int[8] ;
    input \m_cablesIn[8][8] ;
    output \m_cablesIn[9][8] ;
    output \m_cablesIn[9][9] ;
    input \B_int[5] ;
    input \m_cablesIn[8][5] ;
    input \B_int[6] ;
    input \m_cablesIn[8][6] ;
    output \m_cablesIn[9][6] ;
    output \m_cablesIn[9][7] ;
    input \B_int[3] ;
    input \m_cablesIn[8][3] ;
    input \B_int[4] ;
    input \m_cablesIn[8][4] ;
    output \m_cablesIn[9][4] ;
    output \m_cablesIn[9][5] ;
    input \B_int[1] ;
    input \m_cablesIn[8][1] ;
    input \B_int[2] ;
    input \m_cablesIn[8][2] ;
    output \m_cablesIn[9][2] ;
    output \m_cablesIn[9][3] ;
    input \B_int[0] ;
    input \frac_div[19] ;
    output \m_cablesIn[9][1] ;
    
    
    wire n62425, n62424, n62423, n62422, n62421, n62420, n62419, 
        n62418, n62417, n62416, n62415, n62414;
    
    CCU2D add_3303_25 (.A0(\m_cablesIn[8][23] ), .B0(\QQ_in[8][7] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[8][24] ), .B1(\QQ_in[8][7] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62425), .S0(\m_cablesIn[9][24] ), 
          .S1(\QQ_in[9][8] ));
    defparam add_3303_25.INIT0 = 16'h5666;
    defparam add_3303_25.INIT1 = 16'h5999;
    defparam add_3303_25.INJECT1_0 = "NO";
    defparam add_3303_25.INJECT1_1 = "NO";
    CCU2D add_3303_23 (.A0(\B_int[21] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][22] ), 
          .D1(GND_net), .CIN(n62424), .COUT(n62425), .S0(\m_cablesIn[9][22] ), 
          .S1(\m_cablesIn[9][23] ));
    defparam add_3303_23.INIT0 = 16'h6969;
    defparam add_3303_23.INIT1 = 16'h6969;
    defparam add_3303_23.INJECT1_0 = "NO";
    defparam add_3303_23.INJECT1_1 = "NO";
    CCU2D add_3303_21 (.A0(\B_int[19] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][20] ), 
          .D1(GND_net), .CIN(n62423), .COUT(n62424), .S0(\m_cablesIn[9][20] ), 
          .S1(\m_cablesIn[9][21] ));
    defparam add_3303_21.INIT0 = 16'h6969;
    defparam add_3303_21.INIT1 = 16'h6969;
    defparam add_3303_21.INJECT1_0 = "NO";
    defparam add_3303_21.INJECT1_1 = "NO";
    CCU2D add_3303_19 (.A0(\B_int[17] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][18] ), 
          .D1(GND_net), .CIN(n62422), .COUT(n62423), .S0(\m_cablesIn[9][18] ), 
          .S1(\m_cablesIn[9][19] ));
    defparam add_3303_19.INIT0 = 16'h6969;
    defparam add_3303_19.INIT1 = 16'h6969;
    defparam add_3303_19.INJECT1_0 = "NO";
    defparam add_3303_19.INJECT1_1 = "NO";
    CCU2D add_3303_17 (.A0(\B_int[15] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][16] ), 
          .D1(GND_net), .CIN(n62421), .COUT(n62422), .S0(\m_cablesIn[9][16] ), 
          .S1(\m_cablesIn[9][17] ));
    defparam add_3303_17.INIT0 = 16'h6969;
    defparam add_3303_17.INIT1 = 16'h6969;
    defparam add_3303_17.INJECT1_0 = "NO";
    defparam add_3303_17.INJECT1_1 = "NO";
    CCU2D add_3303_15 (.A0(\B_int[13] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][14] ), 
          .D1(GND_net), .CIN(n62420), .COUT(n62421), .S0(\m_cablesIn[9][14] ), 
          .S1(\m_cablesIn[9][15] ));
    defparam add_3303_15.INIT0 = 16'h6969;
    defparam add_3303_15.INIT1 = 16'h6969;
    defparam add_3303_15.INJECT1_0 = "NO";
    defparam add_3303_15.INJECT1_1 = "NO";
    CCU2D add_3303_13 (.A0(\B_int[11] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][12] ), 
          .D1(GND_net), .CIN(n62419), .COUT(n62420), .S0(\m_cablesIn[9][12] ), 
          .S1(\m_cablesIn[9][13] ));
    defparam add_3303_13.INIT0 = 16'h6969;
    defparam add_3303_13.INIT1 = 16'h6969;
    defparam add_3303_13.INJECT1_0 = "NO";
    defparam add_3303_13.INJECT1_1 = "NO";
    CCU2D add_3303_11 (.A0(\B_int[9] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][10] ), 
          .D1(GND_net), .CIN(n62418), .COUT(n62419), .S0(\m_cablesIn[9][10] ), 
          .S1(\m_cablesIn[9][11] ));
    defparam add_3303_11.INIT0 = 16'h6969;
    defparam add_3303_11.INIT1 = 16'h6969;
    defparam add_3303_11.INJECT1_0 = "NO";
    defparam add_3303_11.INJECT1_1 = "NO";
    CCU2D add_3303_9 (.A0(\B_int[7] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][8] ), 
          .D1(GND_net), .CIN(n62417), .COUT(n62418), .S0(\m_cablesIn[9][8] ), 
          .S1(\m_cablesIn[9][9] ));
    defparam add_3303_9.INIT0 = 16'h6969;
    defparam add_3303_9.INIT1 = 16'h6969;
    defparam add_3303_9.INJECT1_0 = "NO";
    defparam add_3303_9.INJECT1_1 = "NO";
    CCU2D add_3303_7 (.A0(\B_int[5] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][6] ), 
          .D1(GND_net), .CIN(n62416), .COUT(n62417), .S0(\m_cablesIn[9][6] ), 
          .S1(\m_cablesIn[9][7] ));
    defparam add_3303_7.INIT0 = 16'h6969;
    defparam add_3303_7.INIT1 = 16'h6969;
    defparam add_3303_7.INJECT1_0 = "NO";
    defparam add_3303_7.INJECT1_1 = "NO";
    CCU2D add_3303_5 (.A0(\B_int[3] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][4] ), 
          .D1(GND_net), .CIN(n62415), .COUT(n62416), .S0(\m_cablesIn[9][4] ), 
          .S1(\m_cablesIn[9][5] ));
    defparam add_3303_5.INIT0 = 16'h6969;
    defparam add_3303_5.INIT1 = 16'h6969;
    defparam add_3303_5.INJECT1_0 = "NO";
    defparam add_3303_5.INJECT1_1 = "NO";
    CCU2D add_3303_3 (.A0(\B_int[1] ), .B0(\QQ_in[8][7] ), .C0(\m_cablesIn[8][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[8][7] ), .C1(\m_cablesIn[8][2] ), 
          .D1(GND_net), .CIN(n62414), .COUT(n62415), .S0(\m_cablesIn[9][2] ), 
          .S1(\m_cablesIn[9][3] ));
    defparam add_3303_3.INIT0 = 16'h6969;
    defparam add_3303_3.INIT1 = 16'h6969;
    defparam add_3303_3.INJECT1_0 = "NO";
    defparam add_3303_3.INJECT1_1 = "NO";
    CCU2D add_3303_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[8][7] ), .C1(\frac_div[19] ), .D1(GND_net), 
          .COUT(n62414), .S1(\m_cablesIn[9][1] ));
    defparam add_3303_1.INIT0 = 16'hF000;
    defparam add_3303_1.INIT1 = 16'h6969;
    defparam add_3303_1.INJECT1_0 = "NO";
    defparam add_3303_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U0 
//

module \a_s(24)_U0  (\m_cablesIn[7][23] , \QQ_in[7][6] , GND_net, \m_cablesIn[7][24] , 
            \m_cablesIn[8][24] , \QQ_in[8][7] , \B_int[21] , \m_cablesIn[7][21] , 
            \B_int[22] , \m_cablesIn[7][22] , \m_cablesIn[8][22] , \m_cablesIn[8][23] , 
            \B_int[19] , \m_cablesIn[7][19] , \B_int[20] , \m_cablesIn[7][20] , 
            \m_cablesIn[8][20] , \m_cablesIn[8][21] , \B_int[17] , \m_cablesIn[7][17] , 
            \B_int[18] , \m_cablesIn[7][18] , \m_cablesIn[8][18] , \m_cablesIn[8][19] , 
            \B_int[15] , \m_cablesIn[7][15] , \B_int[16] , \m_cablesIn[7][16] , 
            \m_cablesIn[8][16] , \m_cablesIn[8][17] , \B_int[13] , \m_cablesIn[7][13] , 
            \B_int[14] , \m_cablesIn[7][14] , \m_cablesIn[8][14] , \m_cablesIn[8][15] , 
            \B_int[11] , \m_cablesIn[7][11] , \B_int[12] , \m_cablesIn[7][12] , 
            \m_cablesIn[8][12] , \m_cablesIn[8][13] , \B_int[9] , \m_cablesIn[7][9] , 
            \B_int[10] , \m_cablesIn[7][10] , \m_cablesIn[8][10] , \m_cablesIn[8][11] , 
            \B_int[7] , \m_cablesIn[7][7] , \B_int[8] , \m_cablesIn[7][8] , 
            \m_cablesIn[8][8] , \m_cablesIn[8][9] , \B_int[5] , \m_cablesIn[7][5] , 
            \B_int[6] , \m_cablesIn[7][6] , \m_cablesIn[8][6] , \m_cablesIn[8][7] , 
            \B_int[3] , \m_cablesIn[7][3] , \B_int[4] , \m_cablesIn[7][4] , 
            \m_cablesIn[8][4] , \m_cablesIn[8][5] , \B_int[1] , \m_cablesIn[7][1] , 
            \B_int[2] , \m_cablesIn[7][2] , \m_cablesIn[8][2] , \m_cablesIn[8][3] , 
            \B_int[0] , \frac_div[20] , \m_cablesIn[8][1] );
    input \m_cablesIn[7][23] ;
    input \QQ_in[7][6] ;
    input GND_net;
    input \m_cablesIn[7][24] ;
    output \m_cablesIn[8][24] ;
    output \QQ_in[8][7] ;
    input \B_int[21] ;
    input \m_cablesIn[7][21] ;
    input \B_int[22] ;
    input \m_cablesIn[7][22] ;
    output \m_cablesIn[8][22] ;
    output \m_cablesIn[8][23] ;
    input \B_int[19] ;
    input \m_cablesIn[7][19] ;
    input \B_int[20] ;
    input \m_cablesIn[7][20] ;
    output \m_cablesIn[8][20] ;
    output \m_cablesIn[8][21] ;
    input \B_int[17] ;
    input \m_cablesIn[7][17] ;
    input \B_int[18] ;
    input \m_cablesIn[7][18] ;
    output \m_cablesIn[8][18] ;
    output \m_cablesIn[8][19] ;
    input \B_int[15] ;
    input \m_cablesIn[7][15] ;
    input \B_int[16] ;
    input \m_cablesIn[7][16] ;
    output \m_cablesIn[8][16] ;
    output \m_cablesIn[8][17] ;
    input \B_int[13] ;
    input \m_cablesIn[7][13] ;
    input \B_int[14] ;
    input \m_cablesIn[7][14] ;
    output \m_cablesIn[8][14] ;
    output \m_cablesIn[8][15] ;
    input \B_int[11] ;
    input \m_cablesIn[7][11] ;
    input \B_int[12] ;
    input \m_cablesIn[7][12] ;
    output \m_cablesIn[8][12] ;
    output \m_cablesIn[8][13] ;
    input \B_int[9] ;
    input \m_cablesIn[7][9] ;
    input \B_int[10] ;
    input \m_cablesIn[7][10] ;
    output \m_cablesIn[8][10] ;
    output \m_cablesIn[8][11] ;
    input \B_int[7] ;
    input \m_cablesIn[7][7] ;
    input \B_int[8] ;
    input \m_cablesIn[7][8] ;
    output \m_cablesIn[8][8] ;
    output \m_cablesIn[8][9] ;
    input \B_int[5] ;
    input \m_cablesIn[7][5] ;
    input \B_int[6] ;
    input \m_cablesIn[7][6] ;
    output \m_cablesIn[8][6] ;
    output \m_cablesIn[8][7] ;
    input \B_int[3] ;
    input \m_cablesIn[7][3] ;
    input \B_int[4] ;
    input \m_cablesIn[7][4] ;
    output \m_cablesIn[8][4] ;
    output \m_cablesIn[8][5] ;
    input \B_int[1] ;
    input \m_cablesIn[7][1] ;
    input \B_int[2] ;
    input \m_cablesIn[7][2] ;
    output \m_cablesIn[8][2] ;
    output \m_cablesIn[8][3] ;
    input \B_int[0] ;
    input \frac_div[20] ;
    output \m_cablesIn[8][1] ;
    
    
    wire n62438, n62437, n62436, n62435, n62434, n62433, n62432, 
        n62431, n62430, n62429, n62428, n62427;
    
    CCU2D add_3277_25 (.A0(\m_cablesIn[7][23] ), .B0(\QQ_in[7][6] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[7][24] ), .B1(\QQ_in[7][6] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62438), .S0(\m_cablesIn[8][24] ), 
          .S1(\QQ_in[8][7] ));
    defparam add_3277_25.INIT0 = 16'h5666;
    defparam add_3277_25.INIT1 = 16'h5999;
    defparam add_3277_25.INJECT1_0 = "NO";
    defparam add_3277_25.INJECT1_1 = "NO";
    CCU2D add_3277_23 (.A0(\B_int[21] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][22] ), 
          .D1(GND_net), .CIN(n62437), .COUT(n62438), .S0(\m_cablesIn[8][22] ), 
          .S1(\m_cablesIn[8][23] ));
    defparam add_3277_23.INIT0 = 16'h6969;
    defparam add_3277_23.INIT1 = 16'h6969;
    defparam add_3277_23.INJECT1_0 = "NO";
    defparam add_3277_23.INJECT1_1 = "NO";
    CCU2D add_3277_21 (.A0(\B_int[19] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][20] ), 
          .D1(GND_net), .CIN(n62436), .COUT(n62437), .S0(\m_cablesIn[8][20] ), 
          .S1(\m_cablesIn[8][21] ));
    defparam add_3277_21.INIT0 = 16'h6969;
    defparam add_3277_21.INIT1 = 16'h6969;
    defparam add_3277_21.INJECT1_0 = "NO";
    defparam add_3277_21.INJECT1_1 = "NO";
    CCU2D add_3277_19 (.A0(\B_int[17] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][18] ), 
          .D1(GND_net), .CIN(n62435), .COUT(n62436), .S0(\m_cablesIn[8][18] ), 
          .S1(\m_cablesIn[8][19] ));
    defparam add_3277_19.INIT0 = 16'h6969;
    defparam add_3277_19.INIT1 = 16'h6969;
    defparam add_3277_19.INJECT1_0 = "NO";
    defparam add_3277_19.INJECT1_1 = "NO";
    CCU2D add_3277_17 (.A0(\B_int[15] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][16] ), 
          .D1(GND_net), .CIN(n62434), .COUT(n62435), .S0(\m_cablesIn[8][16] ), 
          .S1(\m_cablesIn[8][17] ));
    defparam add_3277_17.INIT0 = 16'h6969;
    defparam add_3277_17.INIT1 = 16'h6969;
    defparam add_3277_17.INJECT1_0 = "NO";
    defparam add_3277_17.INJECT1_1 = "NO";
    CCU2D add_3277_15 (.A0(\B_int[13] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][14] ), 
          .D1(GND_net), .CIN(n62433), .COUT(n62434), .S0(\m_cablesIn[8][14] ), 
          .S1(\m_cablesIn[8][15] ));
    defparam add_3277_15.INIT0 = 16'h6969;
    defparam add_3277_15.INIT1 = 16'h6969;
    defparam add_3277_15.INJECT1_0 = "NO";
    defparam add_3277_15.INJECT1_1 = "NO";
    CCU2D add_3277_13 (.A0(\B_int[11] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][12] ), 
          .D1(GND_net), .CIN(n62432), .COUT(n62433), .S0(\m_cablesIn[8][12] ), 
          .S1(\m_cablesIn[8][13] ));
    defparam add_3277_13.INIT0 = 16'h6969;
    defparam add_3277_13.INIT1 = 16'h6969;
    defparam add_3277_13.INJECT1_0 = "NO";
    defparam add_3277_13.INJECT1_1 = "NO";
    CCU2D add_3277_11 (.A0(\B_int[9] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][10] ), 
          .D1(GND_net), .CIN(n62431), .COUT(n62432), .S0(\m_cablesIn[8][10] ), 
          .S1(\m_cablesIn[8][11] ));
    defparam add_3277_11.INIT0 = 16'h6969;
    defparam add_3277_11.INIT1 = 16'h6969;
    defparam add_3277_11.INJECT1_0 = "NO";
    defparam add_3277_11.INJECT1_1 = "NO";
    CCU2D add_3277_9 (.A0(\B_int[7] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][8] ), 
          .D1(GND_net), .CIN(n62430), .COUT(n62431), .S0(\m_cablesIn[8][8] ), 
          .S1(\m_cablesIn[8][9] ));
    defparam add_3277_9.INIT0 = 16'h6969;
    defparam add_3277_9.INIT1 = 16'h6969;
    defparam add_3277_9.INJECT1_0 = "NO";
    defparam add_3277_9.INJECT1_1 = "NO";
    CCU2D add_3277_7 (.A0(\B_int[5] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][6] ), 
          .D1(GND_net), .CIN(n62429), .COUT(n62430), .S0(\m_cablesIn[8][6] ), 
          .S1(\m_cablesIn[8][7] ));
    defparam add_3277_7.INIT0 = 16'h6969;
    defparam add_3277_7.INIT1 = 16'h6969;
    defparam add_3277_7.INJECT1_0 = "NO";
    defparam add_3277_7.INJECT1_1 = "NO";
    CCU2D add_3277_5 (.A0(\B_int[3] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][4] ), 
          .D1(GND_net), .CIN(n62428), .COUT(n62429), .S0(\m_cablesIn[8][4] ), 
          .S1(\m_cablesIn[8][5] ));
    defparam add_3277_5.INIT0 = 16'h6969;
    defparam add_3277_5.INIT1 = 16'h6969;
    defparam add_3277_5.INJECT1_0 = "NO";
    defparam add_3277_5.INJECT1_1 = "NO";
    CCU2D add_3277_3 (.A0(\B_int[1] ), .B0(\QQ_in[7][6] ), .C0(\m_cablesIn[7][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[7][6] ), .C1(\m_cablesIn[7][2] ), 
          .D1(GND_net), .CIN(n62427), .COUT(n62428), .S0(\m_cablesIn[8][2] ), 
          .S1(\m_cablesIn[8][3] ));
    defparam add_3277_3.INIT0 = 16'h6969;
    defparam add_3277_3.INIT1 = 16'h6969;
    defparam add_3277_3.INJECT1_0 = "NO";
    defparam add_3277_3.INJECT1_1 = "NO";
    CCU2D add_3277_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[7][6] ), .C1(\frac_div[20] ), .D1(GND_net), 
          .COUT(n62427), .S1(\m_cablesIn[8][1] ));
    defparam add_3277_1.INIT0 = 16'hF000;
    defparam add_3277_1.INIT1 = 16'h6969;
    defparam add_3277_1.INJECT1_0 = "NO";
    defparam add_3277_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U1 
//

module \a_s(24)_U1  (\m_cablesIn[6][23] , \QQ_in[6][5] , GND_net, \m_cablesIn[6][24] , 
            \m_cablesIn[7][24] , \QQ_in[7][6] , \B_int[21] , \m_cablesIn[6][21] , 
            \B_int[22] , \m_cablesIn[6][22] , \m_cablesIn[7][22] , \m_cablesIn[7][23] , 
            \B_int[19] , \m_cablesIn[6][19] , \B_int[20] , \m_cablesIn[6][20] , 
            \m_cablesIn[7][20] , \m_cablesIn[7][21] , \B_int[17] , \m_cablesIn[6][17] , 
            \B_int[18] , \m_cablesIn[6][18] , \m_cablesIn[7][18] , \m_cablesIn[7][19] , 
            \B_int[15] , \m_cablesIn[6][15] , \B_int[16] , \m_cablesIn[6][16] , 
            \m_cablesIn[7][16] , \m_cablesIn[7][17] , \B_int[13] , \m_cablesIn[6][13] , 
            \B_int[14] , \m_cablesIn[6][14] , \m_cablesIn[7][14] , \m_cablesIn[7][15] , 
            \B_int[11] , \m_cablesIn[6][11] , \B_int[12] , \m_cablesIn[6][12] , 
            \m_cablesIn[7][12] , \m_cablesIn[7][13] , \B_int[9] , \m_cablesIn[6][9] , 
            \B_int[10] , \m_cablesIn[6][10] , \m_cablesIn[7][10] , \m_cablesIn[7][11] , 
            \B_int[7] , \m_cablesIn[6][7] , \B_int[8] , \m_cablesIn[6][8] , 
            \m_cablesIn[7][8] , \m_cablesIn[7][9] , \B_int[5] , \m_cablesIn[6][5] , 
            \B_int[6] , \m_cablesIn[6][6] , \m_cablesIn[7][6] , \m_cablesIn[7][7] , 
            \B_int[3] , \m_cablesIn[6][3] , \B_int[4] , \m_cablesIn[6][4] , 
            \m_cablesIn[7][4] , \m_cablesIn[7][5] , \B_int[1] , \m_cablesIn[6][1] , 
            \B_int[2] , \m_cablesIn[6][2] , \m_cablesIn[7][2] , \m_cablesIn[7][3] , 
            \B_int[0] , \frac_div[21] , \m_cablesIn[7][1] );
    input \m_cablesIn[6][23] ;
    input \QQ_in[6][5] ;
    input GND_net;
    input \m_cablesIn[6][24] ;
    output \m_cablesIn[7][24] ;
    output \QQ_in[7][6] ;
    input \B_int[21] ;
    input \m_cablesIn[6][21] ;
    input \B_int[22] ;
    input \m_cablesIn[6][22] ;
    output \m_cablesIn[7][22] ;
    output \m_cablesIn[7][23] ;
    input \B_int[19] ;
    input \m_cablesIn[6][19] ;
    input \B_int[20] ;
    input \m_cablesIn[6][20] ;
    output \m_cablesIn[7][20] ;
    output \m_cablesIn[7][21] ;
    input \B_int[17] ;
    input \m_cablesIn[6][17] ;
    input \B_int[18] ;
    input \m_cablesIn[6][18] ;
    output \m_cablesIn[7][18] ;
    output \m_cablesIn[7][19] ;
    input \B_int[15] ;
    input \m_cablesIn[6][15] ;
    input \B_int[16] ;
    input \m_cablesIn[6][16] ;
    output \m_cablesIn[7][16] ;
    output \m_cablesIn[7][17] ;
    input \B_int[13] ;
    input \m_cablesIn[6][13] ;
    input \B_int[14] ;
    input \m_cablesIn[6][14] ;
    output \m_cablesIn[7][14] ;
    output \m_cablesIn[7][15] ;
    input \B_int[11] ;
    input \m_cablesIn[6][11] ;
    input \B_int[12] ;
    input \m_cablesIn[6][12] ;
    output \m_cablesIn[7][12] ;
    output \m_cablesIn[7][13] ;
    input \B_int[9] ;
    input \m_cablesIn[6][9] ;
    input \B_int[10] ;
    input \m_cablesIn[6][10] ;
    output \m_cablesIn[7][10] ;
    output \m_cablesIn[7][11] ;
    input \B_int[7] ;
    input \m_cablesIn[6][7] ;
    input \B_int[8] ;
    input \m_cablesIn[6][8] ;
    output \m_cablesIn[7][8] ;
    output \m_cablesIn[7][9] ;
    input \B_int[5] ;
    input \m_cablesIn[6][5] ;
    input \B_int[6] ;
    input \m_cablesIn[6][6] ;
    output \m_cablesIn[7][6] ;
    output \m_cablesIn[7][7] ;
    input \B_int[3] ;
    input \m_cablesIn[6][3] ;
    input \B_int[4] ;
    input \m_cablesIn[6][4] ;
    output \m_cablesIn[7][4] ;
    output \m_cablesIn[7][5] ;
    input \B_int[1] ;
    input \m_cablesIn[6][1] ;
    input \B_int[2] ;
    input \m_cablesIn[6][2] ;
    output \m_cablesIn[7][2] ;
    output \m_cablesIn[7][3] ;
    input \B_int[0] ;
    input \frac_div[21] ;
    output \m_cablesIn[7][1] ;
    
    
    wire n62451, n62450, n62449, n62448, n62447, n62446, n62445, 
        n62444, n62443, n62442, n62441, n62440;
    
    CCU2D add_3251_25 (.A0(\m_cablesIn[6][23] ), .B0(\QQ_in[6][5] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[6][24] ), .B1(\QQ_in[6][5] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62451), .S0(\m_cablesIn[7][24] ), 
          .S1(\QQ_in[7][6] ));
    defparam add_3251_25.INIT0 = 16'h5666;
    defparam add_3251_25.INIT1 = 16'h5999;
    defparam add_3251_25.INJECT1_0 = "NO";
    defparam add_3251_25.INJECT1_1 = "NO";
    CCU2D add_3251_23 (.A0(\B_int[21] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][22] ), 
          .D1(GND_net), .CIN(n62450), .COUT(n62451), .S0(\m_cablesIn[7][22] ), 
          .S1(\m_cablesIn[7][23] ));
    defparam add_3251_23.INIT0 = 16'h6969;
    defparam add_3251_23.INIT1 = 16'h6969;
    defparam add_3251_23.INJECT1_0 = "NO";
    defparam add_3251_23.INJECT1_1 = "NO";
    CCU2D add_3251_21 (.A0(\B_int[19] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][20] ), 
          .D1(GND_net), .CIN(n62449), .COUT(n62450), .S0(\m_cablesIn[7][20] ), 
          .S1(\m_cablesIn[7][21] ));
    defparam add_3251_21.INIT0 = 16'h6969;
    defparam add_3251_21.INIT1 = 16'h6969;
    defparam add_3251_21.INJECT1_0 = "NO";
    defparam add_3251_21.INJECT1_1 = "NO";
    CCU2D add_3251_19 (.A0(\B_int[17] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][18] ), 
          .D1(GND_net), .CIN(n62448), .COUT(n62449), .S0(\m_cablesIn[7][18] ), 
          .S1(\m_cablesIn[7][19] ));
    defparam add_3251_19.INIT0 = 16'h6969;
    defparam add_3251_19.INIT1 = 16'h6969;
    defparam add_3251_19.INJECT1_0 = "NO";
    defparam add_3251_19.INJECT1_1 = "NO";
    CCU2D add_3251_17 (.A0(\B_int[15] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][16] ), 
          .D1(GND_net), .CIN(n62447), .COUT(n62448), .S0(\m_cablesIn[7][16] ), 
          .S1(\m_cablesIn[7][17] ));
    defparam add_3251_17.INIT0 = 16'h6969;
    defparam add_3251_17.INIT1 = 16'h6969;
    defparam add_3251_17.INJECT1_0 = "NO";
    defparam add_3251_17.INJECT1_1 = "NO";
    CCU2D add_3251_15 (.A0(\B_int[13] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][14] ), 
          .D1(GND_net), .CIN(n62446), .COUT(n62447), .S0(\m_cablesIn[7][14] ), 
          .S1(\m_cablesIn[7][15] ));
    defparam add_3251_15.INIT0 = 16'h6969;
    defparam add_3251_15.INIT1 = 16'h6969;
    defparam add_3251_15.INJECT1_0 = "NO";
    defparam add_3251_15.INJECT1_1 = "NO";
    CCU2D add_3251_13 (.A0(\B_int[11] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][12] ), 
          .D1(GND_net), .CIN(n62445), .COUT(n62446), .S0(\m_cablesIn[7][12] ), 
          .S1(\m_cablesIn[7][13] ));
    defparam add_3251_13.INIT0 = 16'h6969;
    defparam add_3251_13.INIT1 = 16'h6969;
    defparam add_3251_13.INJECT1_0 = "NO";
    defparam add_3251_13.INJECT1_1 = "NO";
    CCU2D add_3251_11 (.A0(\B_int[9] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][10] ), 
          .D1(GND_net), .CIN(n62444), .COUT(n62445), .S0(\m_cablesIn[7][10] ), 
          .S1(\m_cablesIn[7][11] ));
    defparam add_3251_11.INIT0 = 16'h6969;
    defparam add_3251_11.INIT1 = 16'h6969;
    defparam add_3251_11.INJECT1_0 = "NO";
    defparam add_3251_11.INJECT1_1 = "NO";
    CCU2D add_3251_9 (.A0(\B_int[7] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][8] ), 
          .D1(GND_net), .CIN(n62443), .COUT(n62444), .S0(\m_cablesIn[7][8] ), 
          .S1(\m_cablesIn[7][9] ));
    defparam add_3251_9.INIT0 = 16'h6969;
    defparam add_3251_9.INIT1 = 16'h6969;
    defparam add_3251_9.INJECT1_0 = "NO";
    defparam add_3251_9.INJECT1_1 = "NO";
    CCU2D add_3251_7 (.A0(\B_int[5] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][6] ), 
          .D1(GND_net), .CIN(n62442), .COUT(n62443), .S0(\m_cablesIn[7][6] ), 
          .S1(\m_cablesIn[7][7] ));
    defparam add_3251_7.INIT0 = 16'h6969;
    defparam add_3251_7.INIT1 = 16'h6969;
    defparam add_3251_7.INJECT1_0 = "NO";
    defparam add_3251_7.INJECT1_1 = "NO";
    CCU2D add_3251_5 (.A0(\B_int[3] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][4] ), 
          .D1(GND_net), .CIN(n62441), .COUT(n62442), .S0(\m_cablesIn[7][4] ), 
          .S1(\m_cablesIn[7][5] ));
    defparam add_3251_5.INIT0 = 16'h6969;
    defparam add_3251_5.INIT1 = 16'h6969;
    defparam add_3251_5.INJECT1_0 = "NO";
    defparam add_3251_5.INJECT1_1 = "NO";
    CCU2D add_3251_3 (.A0(\B_int[1] ), .B0(\QQ_in[6][5] ), .C0(\m_cablesIn[6][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[6][5] ), .C1(\m_cablesIn[6][2] ), 
          .D1(GND_net), .CIN(n62440), .COUT(n62441), .S0(\m_cablesIn[7][2] ), 
          .S1(\m_cablesIn[7][3] ));
    defparam add_3251_3.INIT0 = 16'h6969;
    defparam add_3251_3.INIT1 = 16'h6969;
    defparam add_3251_3.INJECT1_0 = "NO";
    defparam add_3251_3.INJECT1_1 = "NO";
    CCU2D add_3251_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[6][5] ), .C1(\frac_div[21] ), .D1(GND_net), 
          .COUT(n62440), .S1(\m_cablesIn[7][1] ));
    defparam add_3251_1.INIT0 = 16'hF000;
    defparam add_3251_1.INIT1 = 16'h6969;
    defparam add_3251_1.INJECT1_0 = "NO";
    defparam add_3251_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U2 
//

module \a_s(24)_U2  (\m_cablesIn[5][23] , \QQ_in[5][4] , GND_net, \m_cablesIn[5][24] , 
            \m_cablesIn[6][24] , \QQ_in[6][5] , \B_int[21] , \m_cablesIn[5][21] , 
            \B_int[22] , \m_cablesIn[5][22] , \m_cablesIn[6][22] , \m_cablesIn[6][23] , 
            \B_int[19] , \m_cablesIn[5][19] , \B_int[20] , \m_cablesIn[5][20] , 
            \m_cablesIn[6][20] , \m_cablesIn[6][21] , \B_int[17] , \m_cablesIn[5][17] , 
            \B_int[18] , \m_cablesIn[5][18] , \m_cablesIn[6][18] , \m_cablesIn[6][19] , 
            \B_int[15] , \m_cablesIn[5][15] , \B_int[16] , \m_cablesIn[5][16] , 
            \m_cablesIn[6][16] , \m_cablesIn[6][17] , \B_int[13] , \m_cablesIn[5][13] , 
            \B_int[14] , \m_cablesIn[5][14] , \m_cablesIn[6][14] , \m_cablesIn[6][15] , 
            \B_int[11] , \m_cablesIn[5][11] , \B_int[12] , \m_cablesIn[5][12] , 
            \m_cablesIn[6][12] , \m_cablesIn[6][13] , \B_int[9] , \m_cablesIn[5][9] , 
            \B_int[10] , \m_cablesIn[5][10] , \m_cablesIn[6][10] , \m_cablesIn[6][11] , 
            \B_int[7] , \m_cablesIn[5][7] , \B_int[8] , \m_cablesIn[5][8] , 
            \m_cablesIn[6][8] , \m_cablesIn[6][9] , \B_int[5] , \m_cablesIn[5][5] , 
            \B_int[6] , \m_cablesIn[5][6] , \m_cablesIn[6][6] , \m_cablesIn[6][7] , 
            \B_int[3] , \m_cablesIn[5][3] , \B_int[4] , \m_cablesIn[5][4] , 
            \m_cablesIn[6][4] , \m_cablesIn[6][5] , \B_int[1] , \m_cablesIn[5][1] , 
            \B_int[2] , \m_cablesIn[5][2] , \m_cablesIn[6][2] , \m_cablesIn[6][3] , 
            \B_int[0] , \frac_div[22] , \m_cablesIn[6][1] );
    input \m_cablesIn[5][23] ;
    input \QQ_in[5][4] ;
    input GND_net;
    input \m_cablesIn[5][24] ;
    output \m_cablesIn[6][24] ;
    output \QQ_in[6][5] ;
    input \B_int[21] ;
    input \m_cablesIn[5][21] ;
    input \B_int[22] ;
    input \m_cablesIn[5][22] ;
    output \m_cablesIn[6][22] ;
    output \m_cablesIn[6][23] ;
    input \B_int[19] ;
    input \m_cablesIn[5][19] ;
    input \B_int[20] ;
    input \m_cablesIn[5][20] ;
    output \m_cablesIn[6][20] ;
    output \m_cablesIn[6][21] ;
    input \B_int[17] ;
    input \m_cablesIn[5][17] ;
    input \B_int[18] ;
    input \m_cablesIn[5][18] ;
    output \m_cablesIn[6][18] ;
    output \m_cablesIn[6][19] ;
    input \B_int[15] ;
    input \m_cablesIn[5][15] ;
    input \B_int[16] ;
    input \m_cablesIn[5][16] ;
    output \m_cablesIn[6][16] ;
    output \m_cablesIn[6][17] ;
    input \B_int[13] ;
    input \m_cablesIn[5][13] ;
    input \B_int[14] ;
    input \m_cablesIn[5][14] ;
    output \m_cablesIn[6][14] ;
    output \m_cablesIn[6][15] ;
    input \B_int[11] ;
    input \m_cablesIn[5][11] ;
    input \B_int[12] ;
    input \m_cablesIn[5][12] ;
    output \m_cablesIn[6][12] ;
    output \m_cablesIn[6][13] ;
    input \B_int[9] ;
    input \m_cablesIn[5][9] ;
    input \B_int[10] ;
    input \m_cablesIn[5][10] ;
    output \m_cablesIn[6][10] ;
    output \m_cablesIn[6][11] ;
    input \B_int[7] ;
    input \m_cablesIn[5][7] ;
    input \B_int[8] ;
    input \m_cablesIn[5][8] ;
    output \m_cablesIn[6][8] ;
    output \m_cablesIn[6][9] ;
    input \B_int[5] ;
    input \m_cablesIn[5][5] ;
    input \B_int[6] ;
    input \m_cablesIn[5][6] ;
    output \m_cablesIn[6][6] ;
    output \m_cablesIn[6][7] ;
    input \B_int[3] ;
    input \m_cablesIn[5][3] ;
    input \B_int[4] ;
    input \m_cablesIn[5][4] ;
    output \m_cablesIn[6][4] ;
    output \m_cablesIn[6][5] ;
    input \B_int[1] ;
    input \m_cablesIn[5][1] ;
    input \B_int[2] ;
    input \m_cablesIn[5][2] ;
    output \m_cablesIn[6][2] ;
    output \m_cablesIn[6][3] ;
    input \B_int[0] ;
    input \frac_div[22] ;
    output \m_cablesIn[6][1] ;
    
    
    wire n62464, n62463, n62462, n62461, n62460, n62459, n62458, 
        n62457, n62456, n62455, n62454, n62453;
    
    CCU2D add_3225_25 (.A0(\m_cablesIn[5][23] ), .B0(\QQ_in[5][4] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[5][24] ), .B1(\QQ_in[5][4] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62464), .S0(\m_cablesIn[6][24] ), 
          .S1(\QQ_in[6][5] ));
    defparam add_3225_25.INIT0 = 16'h5666;
    defparam add_3225_25.INIT1 = 16'h5999;
    defparam add_3225_25.INJECT1_0 = "NO";
    defparam add_3225_25.INJECT1_1 = "NO";
    CCU2D add_3225_23 (.A0(\B_int[21] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][22] ), 
          .D1(GND_net), .CIN(n62463), .COUT(n62464), .S0(\m_cablesIn[6][22] ), 
          .S1(\m_cablesIn[6][23] ));
    defparam add_3225_23.INIT0 = 16'h6969;
    defparam add_3225_23.INIT1 = 16'h6969;
    defparam add_3225_23.INJECT1_0 = "NO";
    defparam add_3225_23.INJECT1_1 = "NO";
    CCU2D add_3225_21 (.A0(\B_int[19] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][20] ), 
          .D1(GND_net), .CIN(n62462), .COUT(n62463), .S0(\m_cablesIn[6][20] ), 
          .S1(\m_cablesIn[6][21] ));
    defparam add_3225_21.INIT0 = 16'h6969;
    defparam add_3225_21.INIT1 = 16'h6969;
    defparam add_3225_21.INJECT1_0 = "NO";
    defparam add_3225_21.INJECT1_1 = "NO";
    CCU2D add_3225_19 (.A0(\B_int[17] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][18] ), 
          .D1(GND_net), .CIN(n62461), .COUT(n62462), .S0(\m_cablesIn[6][18] ), 
          .S1(\m_cablesIn[6][19] ));
    defparam add_3225_19.INIT0 = 16'h6969;
    defparam add_3225_19.INIT1 = 16'h6969;
    defparam add_3225_19.INJECT1_0 = "NO";
    defparam add_3225_19.INJECT1_1 = "NO";
    CCU2D add_3225_17 (.A0(\B_int[15] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][16] ), 
          .D1(GND_net), .CIN(n62460), .COUT(n62461), .S0(\m_cablesIn[6][16] ), 
          .S1(\m_cablesIn[6][17] ));
    defparam add_3225_17.INIT0 = 16'h6969;
    defparam add_3225_17.INIT1 = 16'h6969;
    defparam add_3225_17.INJECT1_0 = "NO";
    defparam add_3225_17.INJECT1_1 = "NO";
    CCU2D add_3225_15 (.A0(\B_int[13] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][14] ), 
          .D1(GND_net), .CIN(n62459), .COUT(n62460), .S0(\m_cablesIn[6][14] ), 
          .S1(\m_cablesIn[6][15] ));
    defparam add_3225_15.INIT0 = 16'h6969;
    defparam add_3225_15.INIT1 = 16'h6969;
    defparam add_3225_15.INJECT1_0 = "NO";
    defparam add_3225_15.INJECT1_1 = "NO";
    CCU2D add_3225_13 (.A0(\B_int[11] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][12] ), 
          .D1(GND_net), .CIN(n62458), .COUT(n62459), .S0(\m_cablesIn[6][12] ), 
          .S1(\m_cablesIn[6][13] ));
    defparam add_3225_13.INIT0 = 16'h6969;
    defparam add_3225_13.INIT1 = 16'h6969;
    defparam add_3225_13.INJECT1_0 = "NO";
    defparam add_3225_13.INJECT1_1 = "NO";
    CCU2D add_3225_11 (.A0(\B_int[9] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][10] ), 
          .D1(GND_net), .CIN(n62457), .COUT(n62458), .S0(\m_cablesIn[6][10] ), 
          .S1(\m_cablesIn[6][11] ));
    defparam add_3225_11.INIT0 = 16'h6969;
    defparam add_3225_11.INIT1 = 16'h6969;
    defparam add_3225_11.INJECT1_0 = "NO";
    defparam add_3225_11.INJECT1_1 = "NO";
    CCU2D add_3225_9 (.A0(\B_int[7] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][8] ), 
          .D1(GND_net), .CIN(n62456), .COUT(n62457), .S0(\m_cablesIn[6][8] ), 
          .S1(\m_cablesIn[6][9] ));
    defparam add_3225_9.INIT0 = 16'h6969;
    defparam add_3225_9.INIT1 = 16'h6969;
    defparam add_3225_9.INJECT1_0 = "NO";
    defparam add_3225_9.INJECT1_1 = "NO";
    CCU2D add_3225_7 (.A0(\B_int[5] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][6] ), 
          .D1(GND_net), .CIN(n62455), .COUT(n62456), .S0(\m_cablesIn[6][6] ), 
          .S1(\m_cablesIn[6][7] ));
    defparam add_3225_7.INIT0 = 16'h6969;
    defparam add_3225_7.INIT1 = 16'h6969;
    defparam add_3225_7.INJECT1_0 = "NO";
    defparam add_3225_7.INJECT1_1 = "NO";
    CCU2D add_3225_5 (.A0(\B_int[3] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][4] ), 
          .D1(GND_net), .CIN(n62454), .COUT(n62455), .S0(\m_cablesIn[6][4] ), 
          .S1(\m_cablesIn[6][5] ));
    defparam add_3225_5.INIT0 = 16'h6969;
    defparam add_3225_5.INIT1 = 16'h6969;
    defparam add_3225_5.INJECT1_0 = "NO";
    defparam add_3225_5.INJECT1_1 = "NO";
    CCU2D add_3225_3 (.A0(\B_int[1] ), .B0(\QQ_in[5][4] ), .C0(\m_cablesIn[5][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[5][4] ), .C1(\m_cablesIn[5][2] ), 
          .D1(GND_net), .CIN(n62453), .COUT(n62454), .S0(\m_cablesIn[6][2] ), 
          .S1(\m_cablesIn[6][3] ));
    defparam add_3225_3.INIT0 = 16'h6969;
    defparam add_3225_3.INIT1 = 16'h6969;
    defparam add_3225_3.INJECT1_0 = "NO";
    defparam add_3225_3.INJECT1_1 = "NO";
    CCU2D add_3225_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[5][4] ), .C1(\frac_div[22] ), .D1(GND_net), 
          .COUT(n62453), .S1(\m_cablesIn[6][1] ));
    defparam add_3225_1.INIT0 = 16'hF000;
    defparam add_3225_1.INIT1 = 16'h6969;
    defparam add_3225_1.INJECT1_0 = "NO";
    defparam add_3225_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U3 
//

module \a_s(24)_U3  (\m_cablesIn[4][23] , \QQ_in[4][3] , GND_net, \m_cablesIn[4][24] , 
            \m_cablesIn[5][24] , \QQ_in[5][4] , \B_int[21] , \m_cablesIn[4][21] , 
            \B_int[22] , \m_cablesIn[4][22] , \m_cablesIn[5][22] , \m_cablesIn[5][23] , 
            \B_int[19] , \m_cablesIn[4][19] , \B_int[20] , \m_cablesIn[4][20] , 
            \m_cablesIn[5][20] , \m_cablesIn[5][21] , \B_int[17] , \m_cablesIn[4][17] , 
            \B_int[18] , \m_cablesIn[4][18] , \m_cablesIn[5][18] , \m_cablesIn[5][19] , 
            \B_int[15] , \m_cablesIn[4][15] , \B_int[16] , \m_cablesIn[4][16] , 
            \m_cablesIn[5][16] , \m_cablesIn[5][17] , \B_int[13] , \m_cablesIn[4][13] , 
            \B_int[14] , \m_cablesIn[4][14] , \m_cablesIn[5][14] , \m_cablesIn[5][15] , 
            \B_int[11] , \m_cablesIn[4][11] , \B_int[12] , \m_cablesIn[4][12] , 
            \m_cablesIn[5][12] , \m_cablesIn[5][13] , \B_int[9] , \m_cablesIn[4][9] , 
            \B_int[10] , \m_cablesIn[4][10] , \m_cablesIn[5][10] , \m_cablesIn[5][11] , 
            \B_int[7] , \m_cablesIn[4][7] , \B_int[8] , \m_cablesIn[4][8] , 
            \m_cablesIn[5][8] , \m_cablesIn[5][9] , \B_int[5] , \m_cablesIn[4][5] , 
            \B_int[6] , \m_cablesIn[4][6] , \m_cablesIn[5][6] , \m_cablesIn[5][7] , 
            \B_int[3] , \m_cablesIn[4][3] , \B_int[4] , \m_cablesIn[4][4] , 
            \m_cablesIn[5][4] , \m_cablesIn[5][5] , \B_int[1] , \m_cablesIn[4][1] , 
            \B_int[2] , \m_cablesIn[4][2] , \m_cablesIn[5][2] , \m_cablesIn[5][3] , 
            \B_int[0] , \frac_div[23] , \m_cablesIn[5][1] );
    input \m_cablesIn[4][23] ;
    input \QQ_in[4][3] ;
    input GND_net;
    input \m_cablesIn[4][24] ;
    output \m_cablesIn[5][24] ;
    output \QQ_in[5][4] ;
    input \B_int[21] ;
    input \m_cablesIn[4][21] ;
    input \B_int[22] ;
    input \m_cablesIn[4][22] ;
    output \m_cablesIn[5][22] ;
    output \m_cablesIn[5][23] ;
    input \B_int[19] ;
    input \m_cablesIn[4][19] ;
    input \B_int[20] ;
    input \m_cablesIn[4][20] ;
    output \m_cablesIn[5][20] ;
    output \m_cablesIn[5][21] ;
    input \B_int[17] ;
    input \m_cablesIn[4][17] ;
    input \B_int[18] ;
    input \m_cablesIn[4][18] ;
    output \m_cablesIn[5][18] ;
    output \m_cablesIn[5][19] ;
    input \B_int[15] ;
    input \m_cablesIn[4][15] ;
    input \B_int[16] ;
    input \m_cablesIn[4][16] ;
    output \m_cablesIn[5][16] ;
    output \m_cablesIn[5][17] ;
    input \B_int[13] ;
    input \m_cablesIn[4][13] ;
    input \B_int[14] ;
    input \m_cablesIn[4][14] ;
    output \m_cablesIn[5][14] ;
    output \m_cablesIn[5][15] ;
    input \B_int[11] ;
    input \m_cablesIn[4][11] ;
    input \B_int[12] ;
    input \m_cablesIn[4][12] ;
    output \m_cablesIn[5][12] ;
    output \m_cablesIn[5][13] ;
    input \B_int[9] ;
    input \m_cablesIn[4][9] ;
    input \B_int[10] ;
    input \m_cablesIn[4][10] ;
    output \m_cablesIn[5][10] ;
    output \m_cablesIn[5][11] ;
    input \B_int[7] ;
    input \m_cablesIn[4][7] ;
    input \B_int[8] ;
    input \m_cablesIn[4][8] ;
    output \m_cablesIn[5][8] ;
    output \m_cablesIn[5][9] ;
    input \B_int[5] ;
    input \m_cablesIn[4][5] ;
    input \B_int[6] ;
    input \m_cablesIn[4][6] ;
    output \m_cablesIn[5][6] ;
    output \m_cablesIn[5][7] ;
    input \B_int[3] ;
    input \m_cablesIn[4][3] ;
    input \B_int[4] ;
    input \m_cablesIn[4][4] ;
    output \m_cablesIn[5][4] ;
    output \m_cablesIn[5][5] ;
    input \B_int[1] ;
    input \m_cablesIn[4][1] ;
    input \B_int[2] ;
    input \m_cablesIn[4][2] ;
    output \m_cablesIn[5][2] ;
    output \m_cablesIn[5][3] ;
    input \B_int[0] ;
    input \frac_div[23] ;
    output \m_cablesIn[5][1] ;
    
    
    wire n62477, n62476, n62475, n62474, n62473, n62472, n62471, 
        n62470, n62469, n62468, n62467, n62466;
    
    CCU2D add_3199_25 (.A0(\m_cablesIn[4][23] ), .B0(\QQ_in[4][3] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[4][24] ), .B1(\QQ_in[4][3] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62477), .S0(\m_cablesIn[5][24] ), 
          .S1(\QQ_in[5][4] ));
    defparam add_3199_25.INIT0 = 16'h5666;
    defparam add_3199_25.INIT1 = 16'h5999;
    defparam add_3199_25.INJECT1_0 = "NO";
    defparam add_3199_25.INJECT1_1 = "NO";
    CCU2D add_3199_23 (.A0(\B_int[21] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][22] ), 
          .D1(GND_net), .CIN(n62476), .COUT(n62477), .S0(\m_cablesIn[5][22] ), 
          .S1(\m_cablesIn[5][23] ));
    defparam add_3199_23.INIT0 = 16'h6969;
    defparam add_3199_23.INIT1 = 16'h6969;
    defparam add_3199_23.INJECT1_0 = "NO";
    defparam add_3199_23.INJECT1_1 = "NO";
    CCU2D add_3199_21 (.A0(\B_int[19] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][20] ), 
          .D1(GND_net), .CIN(n62475), .COUT(n62476), .S0(\m_cablesIn[5][20] ), 
          .S1(\m_cablesIn[5][21] ));
    defparam add_3199_21.INIT0 = 16'h6969;
    defparam add_3199_21.INIT1 = 16'h6969;
    defparam add_3199_21.INJECT1_0 = "NO";
    defparam add_3199_21.INJECT1_1 = "NO";
    CCU2D add_3199_19 (.A0(\B_int[17] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][18] ), 
          .D1(GND_net), .CIN(n62474), .COUT(n62475), .S0(\m_cablesIn[5][18] ), 
          .S1(\m_cablesIn[5][19] ));
    defparam add_3199_19.INIT0 = 16'h6969;
    defparam add_3199_19.INIT1 = 16'h6969;
    defparam add_3199_19.INJECT1_0 = "NO";
    defparam add_3199_19.INJECT1_1 = "NO";
    CCU2D add_3199_17 (.A0(\B_int[15] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][16] ), 
          .D1(GND_net), .CIN(n62473), .COUT(n62474), .S0(\m_cablesIn[5][16] ), 
          .S1(\m_cablesIn[5][17] ));
    defparam add_3199_17.INIT0 = 16'h6969;
    defparam add_3199_17.INIT1 = 16'h6969;
    defparam add_3199_17.INJECT1_0 = "NO";
    defparam add_3199_17.INJECT1_1 = "NO";
    CCU2D add_3199_15 (.A0(\B_int[13] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][14] ), 
          .D1(GND_net), .CIN(n62472), .COUT(n62473), .S0(\m_cablesIn[5][14] ), 
          .S1(\m_cablesIn[5][15] ));
    defparam add_3199_15.INIT0 = 16'h6969;
    defparam add_3199_15.INIT1 = 16'h6969;
    defparam add_3199_15.INJECT1_0 = "NO";
    defparam add_3199_15.INJECT1_1 = "NO";
    CCU2D add_3199_13 (.A0(\B_int[11] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][12] ), 
          .D1(GND_net), .CIN(n62471), .COUT(n62472), .S0(\m_cablesIn[5][12] ), 
          .S1(\m_cablesIn[5][13] ));
    defparam add_3199_13.INIT0 = 16'h6969;
    defparam add_3199_13.INIT1 = 16'h6969;
    defparam add_3199_13.INJECT1_0 = "NO";
    defparam add_3199_13.INJECT1_1 = "NO";
    CCU2D add_3199_11 (.A0(\B_int[9] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][10] ), 
          .D1(GND_net), .CIN(n62470), .COUT(n62471), .S0(\m_cablesIn[5][10] ), 
          .S1(\m_cablesIn[5][11] ));
    defparam add_3199_11.INIT0 = 16'h6969;
    defparam add_3199_11.INIT1 = 16'h6969;
    defparam add_3199_11.INJECT1_0 = "NO";
    defparam add_3199_11.INJECT1_1 = "NO";
    CCU2D add_3199_9 (.A0(\B_int[7] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][8] ), 
          .D1(GND_net), .CIN(n62469), .COUT(n62470), .S0(\m_cablesIn[5][8] ), 
          .S1(\m_cablesIn[5][9] ));
    defparam add_3199_9.INIT0 = 16'h6969;
    defparam add_3199_9.INIT1 = 16'h6969;
    defparam add_3199_9.INJECT1_0 = "NO";
    defparam add_3199_9.INJECT1_1 = "NO";
    CCU2D add_3199_7 (.A0(\B_int[5] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][6] ), 
          .D1(GND_net), .CIN(n62468), .COUT(n62469), .S0(\m_cablesIn[5][6] ), 
          .S1(\m_cablesIn[5][7] ));
    defparam add_3199_7.INIT0 = 16'h6969;
    defparam add_3199_7.INIT1 = 16'h6969;
    defparam add_3199_7.INJECT1_0 = "NO";
    defparam add_3199_7.INJECT1_1 = "NO";
    CCU2D add_3199_5 (.A0(\B_int[3] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][4] ), 
          .D1(GND_net), .CIN(n62467), .COUT(n62468), .S0(\m_cablesIn[5][4] ), 
          .S1(\m_cablesIn[5][5] ));
    defparam add_3199_5.INIT0 = 16'h6969;
    defparam add_3199_5.INIT1 = 16'h6969;
    defparam add_3199_5.INJECT1_0 = "NO";
    defparam add_3199_5.INJECT1_1 = "NO";
    CCU2D add_3199_3 (.A0(\B_int[1] ), .B0(\QQ_in[4][3] ), .C0(\m_cablesIn[4][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[4][3] ), .C1(\m_cablesIn[4][2] ), 
          .D1(GND_net), .CIN(n62466), .COUT(n62467), .S0(\m_cablesIn[5][2] ), 
          .S1(\m_cablesIn[5][3] ));
    defparam add_3199_3.INIT0 = 16'h6969;
    defparam add_3199_3.INIT1 = 16'h6969;
    defparam add_3199_3.INJECT1_0 = "NO";
    defparam add_3199_3.INJECT1_1 = "NO";
    CCU2D add_3199_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[4][3] ), .C1(\frac_div[23] ), .D1(GND_net), 
          .COUT(n62466), .S1(\m_cablesIn[5][1] ));
    defparam add_3199_1.INIT0 = 16'hF000;
    defparam add_3199_1.INIT1 = 16'h6969;
    defparam add_3199_1.INJECT1_0 = "NO";
    defparam add_3199_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U4 
//

module \a_s(24)_U4  (\m_cablesIn[3][23] , \QQ_in[3][2] , GND_net, \m_cablesIn[3][24] , 
            \m_cablesIn[4][24] , \QQ_in[4][3] , \B_int[21] , \m_cablesIn[3][21] , 
            \B_int[22] , \m_cablesIn[3][22] , \m_cablesIn[4][22] , \m_cablesIn[4][23] , 
            \B_int[19] , \m_cablesIn[3][19] , \B_int[20] , \m_cablesIn[3][20] , 
            \m_cablesIn[4][20] , \m_cablesIn[4][21] , \B_int[17] , \m_cablesIn[3][17] , 
            \B_int[18] , \m_cablesIn[3][18] , \m_cablesIn[4][18] , \m_cablesIn[4][19] , 
            \B_int[15] , \m_cablesIn[3][15] , \B_int[16] , \m_cablesIn[3][16] , 
            \m_cablesIn[4][16] , \m_cablesIn[4][17] , \B_int[13] , \m_cablesIn[3][13] , 
            \B_int[14] , \m_cablesIn[3][14] , \m_cablesIn[4][14] , \m_cablesIn[4][15] , 
            \B_int[11] , \m_cablesIn[3][11] , \B_int[12] , \m_cablesIn[3][12] , 
            \m_cablesIn[4][12] , \m_cablesIn[4][13] , \B_int[9] , \m_cablesIn[3][9] , 
            \B_int[10] , \m_cablesIn[3][10] , \m_cablesIn[4][10] , \m_cablesIn[4][11] , 
            \B_int[7] , \m_cablesIn[3][7] , \B_int[8] , \m_cablesIn[3][8] , 
            \m_cablesIn[4][8] , \m_cablesIn[4][9] , \B_int[5] , \m_cablesIn[3][5] , 
            \B_int[6] , \m_cablesIn[3][6] , \m_cablesIn[4][6] , \m_cablesIn[4][7] , 
            \B_int[3] , \m_cablesIn[3][3] , \B_int[4] , \m_cablesIn[3][4] , 
            \m_cablesIn[4][4] , \m_cablesIn[4][5] , \B_int[1] , \m_cablesIn[3][1] , 
            \B_int[2] , \m_cablesIn[3][2] , \m_cablesIn[4][2] , \m_cablesIn[4][3] , 
            \B_int[0] , \frac_div[24] , \m_cablesIn[4][1] );
    input \m_cablesIn[3][23] ;
    input \QQ_in[3][2] ;
    input GND_net;
    input \m_cablesIn[3][24] ;
    output \m_cablesIn[4][24] ;
    output \QQ_in[4][3] ;
    input \B_int[21] ;
    input \m_cablesIn[3][21] ;
    input \B_int[22] ;
    input \m_cablesIn[3][22] ;
    output \m_cablesIn[4][22] ;
    output \m_cablesIn[4][23] ;
    input \B_int[19] ;
    input \m_cablesIn[3][19] ;
    input \B_int[20] ;
    input \m_cablesIn[3][20] ;
    output \m_cablesIn[4][20] ;
    output \m_cablesIn[4][21] ;
    input \B_int[17] ;
    input \m_cablesIn[3][17] ;
    input \B_int[18] ;
    input \m_cablesIn[3][18] ;
    output \m_cablesIn[4][18] ;
    output \m_cablesIn[4][19] ;
    input \B_int[15] ;
    input \m_cablesIn[3][15] ;
    input \B_int[16] ;
    input \m_cablesIn[3][16] ;
    output \m_cablesIn[4][16] ;
    output \m_cablesIn[4][17] ;
    input \B_int[13] ;
    input \m_cablesIn[3][13] ;
    input \B_int[14] ;
    input \m_cablesIn[3][14] ;
    output \m_cablesIn[4][14] ;
    output \m_cablesIn[4][15] ;
    input \B_int[11] ;
    input \m_cablesIn[3][11] ;
    input \B_int[12] ;
    input \m_cablesIn[3][12] ;
    output \m_cablesIn[4][12] ;
    output \m_cablesIn[4][13] ;
    input \B_int[9] ;
    input \m_cablesIn[3][9] ;
    input \B_int[10] ;
    input \m_cablesIn[3][10] ;
    output \m_cablesIn[4][10] ;
    output \m_cablesIn[4][11] ;
    input \B_int[7] ;
    input \m_cablesIn[3][7] ;
    input \B_int[8] ;
    input \m_cablesIn[3][8] ;
    output \m_cablesIn[4][8] ;
    output \m_cablesIn[4][9] ;
    input \B_int[5] ;
    input \m_cablesIn[3][5] ;
    input \B_int[6] ;
    input \m_cablesIn[3][6] ;
    output \m_cablesIn[4][6] ;
    output \m_cablesIn[4][7] ;
    input \B_int[3] ;
    input \m_cablesIn[3][3] ;
    input \B_int[4] ;
    input \m_cablesIn[3][4] ;
    output \m_cablesIn[4][4] ;
    output \m_cablesIn[4][5] ;
    input \B_int[1] ;
    input \m_cablesIn[3][1] ;
    input \B_int[2] ;
    input \m_cablesIn[3][2] ;
    output \m_cablesIn[4][2] ;
    output \m_cablesIn[4][3] ;
    input \B_int[0] ;
    input \frac_div[24] ;
    output \m_cablesIn[4][1] ;
    
    
    wire n62490, n62489, n62488, n62487, n62486, n62485, n62484, 
        n62483, n62482, n62481, n62480, n62479;
    
    CCU2D add_3173_25 (.A0(\m_cablesIn[3][23] ), .B0(\QQ_in[3][2] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[3][24] ), .B1(\QQ_in[3][2] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62490), .S0(\m_cablesIn[4][24] ), 
          .S1(\QQ_in[4][3] ));
    defparam add_3173_25.INIT0 = 16'h5666;
    defparam add_3173_25.INIT1 = 16'h5999;
    defparam add_3173_25.INJECT1_0 = "NO";
    defparam add_3173_25.INJECT1_1 = "NO";
    CCU2D add_3173_23 (.A0(\B_int[21] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][22] ), 
          .D1(GND_net), .CIN(n62489), .COUT(n62490), .S0(\m_cablesIn[4][22] ), 
          .S1(\m_cablesIn[4][23] ));
    defparam add_3173_23.INIT0 = 16'h6969;
    defparam add_3173_23.INIT1 = 16'h6969;
    defparam add_3173_23.INJECT1_0 = "NO";
    defparam add_3173_23.INJECT1_1 = "NO";
    CCU2D add_3173_21 (.A0(\B_int[19] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][20] ), 
          .D1(GND_net), .CIN(n62488), .COUT(n62489), .S0(\m_cablesIn[4][20] ), 
          .S1(\m_cablesIn[4][21] ));
    defparam add_3173_21.INIT0 = 16'h6969;
    defparam add_3173_21.INIT1 = 16'h6969;
    defparam add_3173_21.INJECT1_0 = "NO";
    defparam add_3173_21.INJECT1_1 = "NO";
    CCU2D add_3173_19 (.A0(\B_int[17] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][18] ), 
          .D1(GND_net), .CIN(n62487), .COUT(n62488), .S0(\m_cablesIn[4][18] ), 
          .S1(\m_cablesIn[4][19] ));
    defparam add_3173_19.INIT0 = 16'h6969;
    defparam add_3173_19.INIT1 = 16'h6969;
    defparam add_3173_19.INJECT1_0 = "NO";
    defparam add_3173_19.INJECT1_1 = "NO";
    CCU2D add_3173_17 (.A0(\B_int[15] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][16] ), 
          .D1(GND_net), .CIN(n62486), .COUT(n62487), .S0(\m_cablesIn[4][16] ), 
          .S1(\m_cablesIn[4][17] ));
    defparam add_3173_17.INIT0 = 16'h6969;
    defparam add_3173_17.INIT1 = 16'h6969;
    defparam add_3173_17.INJECT1_0 = "NO";
    defparam add_3173_17.INJECT1_1 = "NO";
    CCU2D add_3173_15 (.A0(\B_int[13] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][14] ), 
          .D1(GND_net), .CIN(n62485), .COUT(n62486), .S0(\m_cablesIn[4][14] ), 
          .S1(\m_cablesIn[4][15] ));
    defparam add_3173_15.INIT0 = 16'h6969;
    defparam add_3173_15.INIT1 = 16'h6969;
    defparam add_3173_15.INJECT1_0 = "NO";
    defparam add_3173_15.INJECT1_1 = "NO";
    CCU2D add_3173_13 (.A0(\B_int[11] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][12] ), 
          .D1(GND_net), .CIN(n62484), .COUT(n62485), .S0(\m_cablesIn[4][12] ), 
          .S1(\m_cablesIn[4][13] ));
    defparam add_3173_13.INIT0 = 16'h6969;
    defparam add_3173_13.INIT1 = 16'h6969;
    defparam add_3173_13.INJECT1_0 = "NO";
    defparam add_3173_13.INJECT1_1 = "NO";
    CCU2D add_3173_11 (.A0(\B_int[9] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][10] ), 
          .D1(GND_net), .CIN(n62483), .COUT(n62484), .S0(\m_cablesIn[4][10] ), 
          .S1(\m_cablesIn[4][11] ));
    defparam add_3173_11.INIT0 = 16'h6969;
    defparam add_3173_11.INIT1 = 16'h6969;
    defparam add_3173_11.INJECT1_0 = "NO";
    defparam add_3173_11.INJECT1_1 = "NO";
    CCU2D add_3173_9 (.A0(\B_int[7] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][8] ), 
          .D1(GND_net), .CIN(n62482), .COUT(n62483), .S0(\m_cablesIn[4][8] ), 
          .S1(\m_cablesIn[4][9] ));
    defparam add_3173_9.INIT0 = 16'h6969;
    defparam add_3173_9.INIT1 = 16'h6969;
    defparam add_3173_9.INJECT1_0 = "NO";
    defparam add_3173_9.INJECT1_1 = "NO";
    CCU2D add_3173_7 (.A0(\B_int[5] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][6] ), 
          .D1(GND_net), .CIN(n62481), .COUT(n62482), .S0(\m_cablesIn[4][6] ), 
          .S1(\m_cablesIn[4][7] ));
    defparam add_3173_7.INIT0 = 16'h6969;
    defparam add_3173_7.INIT1 = 16'h6969;
    defparam add_3173_7.INJECT1_0 = "NO";
    defparam add_3173_7.INJECT1_1 = "NO";
    CCU2D add_3173_5 (.A0(\B_int[3] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][4] ), 
          .D1(GND_net), .CIN(n62480), .COUT(n62481), .S0(\m_cablesIn[4][4] ), 
          .S1(\m_cablesIn[4][5] ));
    defparam add_3173_5.INIT0 = 16'h6969;
    defparam add_3173_5.INIT1 = 16'h6969;
    defparam add_3173_5.INJECT1_0 = "NO";
    defparam add_3173_5.INJECT1_1 = "NO";
    CCU2D add_3173_3 (.A0(\B_int[1] ), .B0(\QQ_in[3][2] ), .C0(\m_cablesIn[3][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[3][2] ), .C1(\m_cablesIn[3][2] ), 
          .D1(GND_net), .CIN(n62479), .COUT(n62480), .S0(\m_cablesIn[4][2] ), 
          .S1(\m_cablesIn[4][3] ));
    defparam add_3173_3.INIT0 = 16'h6969;
    defparam add_3173_3.INIT1 = 16'h6969;
    defparam add_3173_3.INJECT1_0 = "NO";
    defparam add_3173_3.INJECT1_1 = "NO";
    CCU2D add_3173_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[3][2] ), .C1(\frac_div[24] ), .D1(GND_net), 
          .COUT(n62479), .S1(\m_cablesIn[4][1] ));
    defparam add_3173_1.INIT0 = 16'hF000;
    defparam add_3173_1.INIT1 = 16'h6969;
    defparam add_3173_1.INJECT1_0 = "NO";
    defparam add_3173_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U5 
//

module \a_s(24)_U5  (\m_cablesIn[2][23] , \QQ_in[2][1] , GND_net, \m_cablesIn[2][24] , 
            \m_cablesIn[3][24] , \QQ_in[3][2] , \B_int[21] , \m_cablesIn[2][21] , 
            \B_int[22] , \m_cablesIn[2][22] , \m_cablesIn[3][22] , \m_cablesIn[3][23] , 
            \B_int[19] , \m_cablesIn[2][19] , \B_int[20] , \m_cablesIn[2][20] , 
            \m_cablesIn[3][20] , \m_cablesIn[3][21] , \B_int[17] , \m_cablesIn[2][17] , 
            \B_int[18] , \m_cablesIn[2][18] , \m_cablesIn[3][18] , \m_cablesIn[3][19] , 
            \B_int[15] , \m_cablesIn[2][15] , \B_int[16] , \m_cablesIn[2][16] , 
            \m_cablesIn[3][16] , \m_cablesIn[3][17] , \B_int[13] , \m_cablesIn[2][13] , 
            \B_int[14] , \m_cablesIn[2][14] , \m_cablesIn[3][14] , \m_cablesIn[3][15] , 
            \B_int[11] , \m_cablesIn[2][11] , \B_int[12] , \m_cablesIn[2][12] , 
            \m_cablesIn[3][12] , \m_cablesIn[3][13] , \B_int[9] , \m_cablesIn[2][9] , 
            \B_int[10] , \m_cablesIn[2][10] , \m_cablesIn[3][10] , \m_cablesIn[3][11] , 
            \B_int[7] , \m_cablesIn[2][7] , \B_int[8] , \m_cablesIn[2][8] , 
            \m_cablesIn[3][8] , \m_cablesIn[3][9] , \B_int[5] , \m_cablesIn[2][5] , 
            \B_int[6] , \m_cablesIn[2][6] , \m_cablesIn[3][6] , \m_cablesIn[3][7] , 
            \B_int[3] , \m_cablesIn[2][3] , \B_int[4] , \m_cablesIn[2][4] , 
            \m_cablesIn[3][4] , \m_cablesIn[3][5] , \B_int[1] , \m_cablesIn[2][1] , 
            \B_int[2] , \m_cablesIn[2][2] , \m_cablesIn[3][2] , \m_cablesIn[3][3] , 
            \B_int[0] , \frac_div[25] , \m_cablesIn[3][1] );
    input \m_cablesIn[2][23] ;
    input \QQ_in[2][1] ;
    input GND_net;
    input \m_cablesIn[2][24] ;
    output \m_cablesIn[3][24] ;
    output \QQ_in[3][2] ;
    input \B_int[21] ;
    input \m_cablesIn[2][21] ;
    input \B_int[22] ;
    input \m_cablesIn[2][22] ;
    output \m_cablesIn[3][22] ;
    output \m_cablesIn[3][23] ;
    input \B_int[19] ;
    input \m_cablesIn[2][19] ;
    input \B_int[20] ;
    input \m_cablesIn[2][20] ;
    output \m_cablesIn[3][20] ;
    output \m_cablesIn[3][21] ;
    input \B_int[17] ;
    input \m_cablesIn[2][17] ;
    input \B_int[18] ;
    input \m_cablesIn[2][18] ;
    output \m_cablesIn[3][18] ;
    output \m_cablesIn[3][19] ;
    input \B_int[15] ;
    input \m_cablesIn[2][15] ;
    input \B_int[16] ;
    input \m_cablesIn[2][16] ;
    output \m_cablesIn[3][16] ;
    output \m_cablesIn[3][17] ;
    input \B_int[13] ;
    input \m_cablesIn[2][13] ;
    input \B_int[14] ;
    input \m_cablesIn[2][14] ;
    output \m_cablesIn[3][14] ;
    output \m_cablesIn[3][15] ;
    input \B_int[11] ;
    input \m_cablesIn[2][11] ;
    input \B_int[12] ;
    input \m_cablesIn[2][12] ;
    output \m_cablesIn[3][12] ;
    output \m_cablesIn[3][13] ;
    input \B_int[9] ;
    input \m_cablesIn[2][9] ;
    input \B_int[10] ;
    input \m_cablesIn[2][10] ;
    output \m_cablesIn[3][10] ;
    output \m_cablesIn[3][11] ;
    input \B_int[7] ;
    input \m_cablesIn[2][7] ;
    input \B_int[8] ;
    input \m_cablesIn[2][8] ;
    output \m_cablesIn[3][8] ;
    output \m_cablesIn[3][9] ;
    input \B_int[5] ;
    input \m_cablesIn[2][5] ;
    input \B_int[6] ;
    input \m_cablesIn[2][6] ;
    output \m_cablesIn[3][6] ;
    output \m_cablesIn[3][7] ;
    input \B_int[3] ;
    input \m_cablesIn[2][3] ;
    input \B_int[4] ;
    input \m_cablesIn[2][4] ;
    output \m_cablesIn[3][4] ;
    output \m_cablesIn[3][5] ;
    input \B_int[1] ;
    input \m_cablesIn[2][1] ;
    input \B_int[2] ;
    input \m_cablesIn[2][2] ;
    output \m_cablesIn[3][2] ;
    output \m_cablesIn[3][3] ;
    input \B_int[0] ;
    input \frac_div[25] ;
    output \m_cablesIn[3][1] ;
    
    
    wire n62503, n62502, n62501, n62500, n62499, n62498, n62497, 
        n62496, n62495, n62494, n62493, n62492;
    
    CCU2D add_3147_25 (.A0(\m_cablesIn[2][23] ), .B0(\QQ_in[2][1] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[2][24] ), .B1(\QQ_in[2][1] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62503), .S0(\m_cablesIn[3][24] ), 
          .S1(\QQ_in[3][2] ));
    defparam add_3147_25.INIT0 = 16'h5666;
    defparam add_3147_25.INIT1 = 16'h5999;
    defparam add_3147_25.INJECT1_0 = "NO";
    defparam add_3147_25.INJECT1_1 = "NO";
    CCU2D add_3147_23 (.A0(\B_int[21] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][22] ), 
          .D1(GND_net), .CIN(n62502), .COUT(n62503), .S0(\m_cablesIn[3][22] ), 
          .S1(\m_cablesIn[3][23] ));
    defparam add_3147_23.INIT0 = 16'h6969;
    defparam add_3147_23.INIT1 = 16'h6969;
    defparam add_3147_23.INJECT1_0 = "NO";
    defparam add_3147_23.INJECT1_1 = "NO";
    CCU2D add_3147_21 (.A0(\B_int[19] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][20] ), 
          .D1(GND_net), .CIN(n62501), .COUT(n62502), .S0(\m_cablesIn[3][20] ), 
          .S1(\m_cablesIn[3][21] ));
    defparam add_3147_21.INIT0 = 16'h6969;
    defparam add_3147_21.INIT1 = 16'h6969;
    defparam add_3147_21.INJECT1_0 = "NO";
    defparam add_3147_21.INJECT1_1 = "NO";
    CCU2D add_3147_19 (.A0(\B_int[17] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][18] ), 
          .D1(GND_net), .CIN(n62500), .COUT(n62501), .S0(\m_cablesIn[3][18] ), 
          .S1(\m_cablesIn[3][19] ));
    defparam add_3147_19.INIT0 = 16'h6969;
    defparam add_3147_19.INIT1 = 16'h6969;
    defparam add_3147_19.INJECT1_0 = "NO";
    defparam add_3147_19.INJECT1_1 = "NO";
    CCU2D add_3147_17 (.A0(\B_int[15] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][16] ), 
          .D1(GND_net), .CIN(n62499), .COUT(n62500), .S0(\m_cablesIn[3][16] ), 
          .S1(\m_cablesIn[3][17] ));
    defparam add_3147_17.INIT0 = 16'h6969;
    defparam add_3147_17.INIT1 = 16'h6969;
    defparam add_3147_17.INJECT1_0 = "NO";
    defparam add_3147_17.INJECT1_1 = "NO";
    CCU2D add_3147_15 (.A0(\B_int[13] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][14] ), 
          .D1(GND_net), .CIN(n62498), .COUT(n62499), .S0(\m_cablesIn[3][14] ), 
          .S1(\m_cablesIn[3][15] ));
    defparam add_3147_15.INIT0 = 16'h6969;
    defparam add_3147_15.INIT1 = 16'h6969;
    defparam add_3147_15.INJECT1_0 = "NO";
    defparam add_3147_15.INJECT1_1 = "NO";
    CCU2D add_3147_13 (.A0(\B_int[11] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][12] ), 
          .D1(GND_net), .CIN(n62497), .COUT(n62498), .S0(\m_cablesIn[3][12] ), 
          .S1(\m_cablesIn[3][13] ));
    defparam add_3147_13.INIT0 = 16'h6969;
    defparam add_3147_13.INIT1 = 16'h6969;
    defparam add_3147_13.INJECT1_0 = "NO";
    defparam add_3147_13.INJECT1_1 = "NO";
    CCU2D add_3147_11 (.A0(\B_int[9] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][10] ), 
          .D1(GND_net), .CIN(n62496), .COUT(n62497), .S0(\m_cablesIn[3][10] ), 
          .S1(\m_cablesIn[3][11] ));
    defparam add_3147_11.INIT0 = 16'h6969;
    defparam add_3147_11.INIT1 = 16'h6969;
    defparam add_3147_11.INJECT1_0 = "NO";
    defparam add_3147_11.INJECT1_1 = "NO";
    CCU2D add_3147_9 (.A0(\B_int[7] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][8] ), 
          .D1(GND_net), .CIN(n62495), .COUT(n62496), .S0(\m_cablesIn[3][8] ), 
          .S1(\m_cablesIn[3][9] ));
    defparam add_3147_9.INIT0 = 16'h6969;
    defparam add_3147_9.INIT1 = 16'h6969;
    defparam add_3147_9.INJECT1_0 = "NO";
    defparam add_3147_9.INJECT1_1 = "NO";
    CCU2D add_3147_7 (.A0(\B_int[5] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][6] ), 
          .D1(GND_net), .CIN(n62494), .COUT(n62495), .S0(\m_cablesIn[3][6] ), 
          .S1(\m_cablesIn[3][7] ));
    defparam add_3147_7.INIT0 = 16'h6969;
    defparam add_3147_7.INIT1 = 16'h6969;
    defparam add_3147_7.INJECT1_0 = "NO";
    defparam add_3147_7.INJECT1_1 = "NO";
    CCU2D add_3147_5 (.A0(\B_int[3] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][4] ), 
          .D1(GND_net), .CIN(n62493), .COUT(n62494), .S0(\m_cablesIn[3][4] ), 
          .S1(\m_cablesIn[3][5] ));
    defparam add_3147_5.INIT0 = 16'h6969;
    defparam add_3147_5.INIT1 = 16'h6969;
    defparam add_3147_5.INJECT1_0 = "NO";
    defparam add_3147_5.INJECT1_1 = "NO";
    CCU2D add_3147_3 (.A0(\B_int[1] ), .B0(\QQ_in[2][1] ), .C0(\m_cablesIn[2][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[2][1] ), .C1(\m_cablesIn[2][2] ), 
          .D1(GND_net), .CIN(n62492), .COUT(n62493), .S0(\m_cablesIn[3][2] ), 
          .S1(\m_cablesIn[3][3] ));
    defparam add_3147_3.INIT0 = 16'h6969;
    defparam add_3147_3.INIT1 = 16'h6969;
    defparam add_3147_3.INJECT1_0 = "NO";
    defparam add_3147_3.INJECT1_1 = "NO";
    CCU2D add_3147_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[2][1] ), .C1(\frac_div[25] ), .D1(GND_net), 
          .COUT(n62492), .S1(\m_cablesIn[3][1] ));
    defparam add_3147_1.INIT0 = 16'hF000;
    defparam add_3147_1.INIT1 = 16'h6969;
    defparam add_3147_1.INJECT1_0 = "NO";
    defparam add_3147_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U6 
//

module \a_s(24)_U6  (\m_cablesIn[1][23] , \QQ_in[1][0] , GND_net, \m_cablesIn[1][24] , 
            \m_cablesIn[2][24] , \QQ_in[2][1] , \B_int[21] , \m_cablesIn[1][21] , 
            \B_int[22] , \m_cablesIn[1][22] , \m_cablesIn[2][22] , \m_cablesIn[2][23] , 
            \B_int[19] , \m_cablesIn[1][19] , \B_int[20] , \m_cablesIn[1][20] , 
            \m_cablesIn[2][20] , \m_cablesIn[2][21] , \B_int[17] , \m_cablesIn[1][17] , 
            \B_int[18] , \m_cablesIn[1][18] , \m_cablesIn[2][18] , \m_cablesIn[2][19] , 
            \B_int[15] , \m_cablesIn[1][15] , \B_int[16] , \m_cablesIn[1][16] , 
            \m_cablesIn[2][16] , \m_cablesIn[2][17] , \B_int[13] , \m_cablesIn[1][13] , 
            \B_int[14] , \m_cablesIn[1][14] , \m_cablesIn[2][14] , \m_cablesIn[2][15] , 
            \B_int[11] , \m_cablesIn[1][11] , \B_int[12] , \m_cablesIn[1][12] , 
            \m_cablesIn[2][12] , \m_cablesIn[2][13] , \B_int[9] , \m_cablesIn[1][9] , 
            \B_int[10] , \m_cablesIn[1][10] , \m_cablesIn[2][10] , \m_cablesIn[2][11] , 
            \B_int[7] , \m_cablesIn[1][7] , \B_int[8] , \m_cablesIn[1][8] , 
            \m_cablesIn[2][8] , \m_cablesIn[2][9] , \B_int[5] , \m_cablesIn[1][5] , 
            \B_int[6] , \m_cablesIn[1][6] , \m_cablesIn[2][6] , \m_cablesIn[2][7] , 
            \B_int[3] , \m_cablesIn[1][3] , \B_int[4] , \m_cablesIn[1][4] , 
            \m_cablesIn[2][4] , \m_cablesIn[2][5] , \B_int[1] , \m_cablesIn[1][1] , 
            \B_int[2] , \m_cablesIn[1][2] , \m_cablesIn[2][2] , \m_cablesIn[2][3] , 
            \B_int[0] , n9256, \m_cablesIn[2][1] );
    input \m_cablesIn[1][23] ;
    input \QQ_in[1][0] ;
    input GND_net;
    input \m_cablesIn[1][24] ;
    output \m_cablesIn[2][24] ;
    output \QQ_in[2][1] ;
    input \B_int[21] ;
    input \m_cablesIn[1][21] ;
    input \B_int[22] ;
    input \m_cablesIn[1][22] ;
    output \m_cablesIn[2][22] ;
    output \m_cablesIn[2][23] ;
    input \B_int[19] ;
    input \m_cablesIn[1][19] ;
    input \B_int[20] ;
    input \m_cablesIn[1][20] ;
    output \m_cablesIn[2][20] ;
    output \m_cablesIn[2][21] ;
    input \B_int[17] ;
    input \m_cablesIn[1][17] ;
    input \B_int[18] ;
    input \m_cablesIn[1][18] ;
    output \m_cablesIn[2][18] ;
    output \m_cablesIn[2][19] ;
    input \B_int[15] ;
    input \m_cablesIn[1][15] ;
    input \B_int[16] ;
    input \m_cablesIn[1][16] ;
    output \m_cablesIn[2][16] ;
    output \m_cablesIn[2][17] ;
    input \B_int[13] ;
    input \m_cablesIn[1][13] ;
    input \B_int[14] ;
    input \m_cablesIn[1][14] ;
    output \m_cablesIn[2][14] ;
    output \m_cablesIn[2][15] ;
    input \B_int[11] ;
    input \m_cablesIn[1][11] ;
    input \B_int[12] ;
    input \m_cablesIn[1][12] ;
    output \m_cablesIn[2][12] ;
    output \m_cablesIn[2][13] ;
    input \B_int[9] ;
    input \m_cablesIn[1][9] ;
    input \B_int[10] ;
    input \m_cablesIn[1][10] ;
    output \m_cablesIn[2][10] ;
    output \m_cablesIn[2][11] ;
    input \B_int[7] ;
    input \m_cablesIn[1][7] ;
    input \B_int[8] ;
    input \m_cablesIn[1][8] ;
    output \m_cablesIn[2][8] ;
    output \m_cablesIn[2][9] ;
    input \B_int[5] ;
    input \m_cablesIn[1][5] ;
    input \B_int[6] ;
    input \m_cablesIn[1][6] ;
    output \m_cablesIn[2][6] ;
    output \m_cablesIn[2][7] ;
    input \B_int[3] ;
    input \m_cablesIn[1][3] ;
    input \B_int[4] ;
    input \m_cablesIn[1][4] ;
    output \m_cablesIn[2][4] ;
    output \m_cablesIn[2][5] ;
    input \B_int[1] ;
    input \m_cablesIn[1][1] ;
    input \B_int[2] ;
    input \m_cablesIn[1][2] ;
    output \m_cablesIn[2][2] ;
    output \m_cablesIn[2][3] ;
    input \B_int[0] ;
    input n9256;
    output \m_cablesIn[2][1] ;
    
    
    wire n62516, n62515, n62514, n62513, n62512, n62511, n62510, 
        n62509, n62508, n62507, n62506, n62505;
    
    CCU2D add_3063_25 (.A0(\m_cablesIn[1][23] ), .B0(\QQ_in[1][0] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[1][24] ), .B1(\QQ_in[1][0] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62516), .S0(\m_cablesIn[2][24] ), 
          .S1(\QQ_in[2][1] ));
    defparam add_3063_25.INIT0 = 16'h5666;
    defparam add_3063_25.INIT1 = 16'h5999;
    defparam add_3063_25.INJECT1_0 = "NO";
    defparam add_3063_25.INJECT1_1 = "NO";
    CCU2D add_3063_23 (.A0(\B_int[21] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][22] ), 
          .D1(GND_net), .CIN(n62515), .COUT(n62516), .S0(\m_cablesIn[2][22] ), 
          .S1(\m_cablesIn[2][23] ));
    defparam add_3063_23.INIT0 = 16'h6969;
    defparam add_3063_23.INIT1 = 16'h6969;
    defparam add_3063_23.INJECT1_0 = "NO";
    defparam add_3063_23.INJECT1_1 = "NO";
    CCU2D add_3063_21 (.A0(\B_int[19] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][20] ), 
          .D1(GND_net), .CIN(n62514), .COUT(n62515), .S0(\m_cablesIn[2][20] ), 
          .S1(\m_cablesIn[2][21] ));
    defparam add_3063_21.INIT0 = 16'h6969;
    defparam add_3063_21.INIT1 = 16'h6969;
    defparam add_3063_21.INJECT1_0 = "NO";
    defparam add_3063_21.INJECT1_1 = "NO";
    CCU2D add_3063_19 (.A0(\B_int[17] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][18] ), 
          .D1(GND_net), .CIN(n62513), .COUT(n62514), .S0(\m_cablesIn[2][18] ), 
          .S1(\m_cablesIn[2][19] ));
    defparam add_3063_19.INIT0 = 16'h6969;
    defparam add_3063_19.INIT1 = 16'h6969;
    defparam add_3063_19.INJECT1_0 = "NO";
    defparam add_3063_19.INJECT1_1 = "NO";
    CCU2D add_3063_17 (.A0(\B_int[15] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][16] ), 
          .D1(GND_net), .CIN(n62512), .COUT(n62513), .S0(\m_cablesIn[2][16] ), 
          .S1(\m_cablesIn[2][17] ));
    defparam add_3063_17.INIT0 = 16'h6969;
    defparam add_3063_17.INIT1 = 16'h6969;
    defparam add_3063_17.INJECT1_0 = "NO";
    defparam add_3063_17.INJECT1_1 = "NO";
    CCU2D add_3063_15 (.A0(\B_int[13] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][14] ), 
          .D1(GND_net), .CIN(n62511), .COUT(n62512), .S0(\m_cablesIn[2][14] ), 
          .S1(\m_cablesIn[2][15] ));
    defparam add_3063_15.INIT0 = 16'h6969;
    defparam add_3063_15.INIT1 = 16'h6969;
    defparam add_3063_15.INJECT1_0 = "NO";
    defparam add_3063_15.INJECT1_1 = "NO";
    CCU2D add_3063_13 (.A0(\B_int[11] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][12] ), 
          .D1(GND_net), .CIN(n62510), .COUT(n62511), .S0(\m_cablesIn[2][12] ), 
          .S1(\m_cablesIn[2][13] ));
    defparam add_3063_13.INIT0 = 16'h6969;
    defparam add_3063_13.INIT1 = 16'h6969;
    defparam add_3063_13.INJECT1_0 = "NO";
    defparam add_3063_13.INJECT1_1 = "NO";
    CCU2D add_3063_11 (.A0(\B_int[9] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][10] ), 
          .D1(GND_net), .CIN(n62509), .COUT(n62510), .S0(\m_cablesIn[2][10] ), 
          .S1(\m_cablesIn[2][11] ));
    defparam add_3063_11.INIT0 = 16'h6969;
    defparam add_3063_11.INIT1 = 16'h6969;
    defparam add_3063_11.INJECT1_0 = "NO";
    defparam add_3063_11.INJECT1_1 = "NO";
    CCU2D add_3063_9 (.A0(\B_int[7] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][8] ), 
          .D1(GND_net), .CIN(n62508), .COUT(n62509), .S0(\m_cablesIn[2][8] ), 
          .S1(\m_cablesIn[2][9] ));
    defparam add_3063_9.INIT0 = 16'h6969;
    defparam add_3063_9.INIT1 = 16'h6969;
    defparam add_3063_9.INJECT1_0 = "NO";
    defparam add_3063_9.INJECT1_1 = "NO";
    CCU2D add_3063_7 (.A0(\B_int[5] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][6] ), 
          .D1(GND_net), .CIN(n62507), .COUT(n62508), .S0(\m_cablesIn[2][6] ), 
          .S1(\m_cablesIn[2][7] ));
    defparam add_3063_7.INIT0 = 16'h6969;
    defparam add_3063_7.INIT1 = 16'h6969;
    defparam add_3063_7.INJECT1_0 = "NO";
    defparam add_3063_7.INJECT1_1 = "NO";
    CCU2D add_3063_5 (.A0(\B_int[3] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][4] ), 
          .D1(GND_net), .CIN(n62506), .COUT(n62507), .S0(\m_cablesIn[2][4] ), 
          .S1(\m_cablesIn[2][5] ));
    defparam add_3063_5.INIT0 = 16'h6969;
    defparam add_3063_5.INIT1 = 16'h6969;
    defparam add_3063_5.INJECT1_0 = "NO";
    defparam add_3063_5.INJECT1_1 = "NO";
    CCU2D add_3063_3 (.A0(\B_int[1] ), .B0(\QQ_in[1][0] ), .C0(\m_cablesIn[1][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[1][0] ), .C1(\m_cablesIn[1][2] ), 
          .D1(GND_net), .CIN(n62505), .COUT(n62506), .S0(\m_cablesIn[2][2] ), 
          .S1(\m_cablesIn[2][3] ));
    defparam add_3063_3.INIT0 = 16'h6969;
    defparam add_3063_3.INIT1 = 16'h6969;
    defparam add_3063_3.INJECT1_0 = "NO";
    defparam add_3063_3.INJECT1_1 = "NO";
    CCU2D add_3063_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[1][0] ), .C1(n9256), .D1(GND_net), 
          .COUT(n62505), .S1(\m_cablesIn[2][1] ));
    defparam add_3063_1.INIT0 = 16'hF000;
    defparam add_3063_1.INIT1 = 16'h6969;
    defparam add_3063_1.INJECT1_0 = "NO";
    defparam add_3063_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U7 
//

module \a_s(24)_U7  (\m_cablesIn[25][23] , \QQ_in[25][24] , GND_net, \m_cablesIn[25][24] , 
            \QQ_in[26][25] , \B_int[21] , \m_cablesIn[25][21] , \B_int[22] , 
            \m_cablesIn[25][22] , \B_int[19] , \m_cablesIn[25][19] , \B_int[20] , 
            \m_cablesIn[25][20] , \B_int[17] , \m_cablesIn[25][17] , \B_int[18] , 
            \m_cablesIn[25][18] , \B_int[15] , \m_cablesIn[25][15] , \B_int[16] , 
            \m_cablesIn[25][16] , \B_int[13] , \m_cablesIn[25][13] , \B_int[14] , 
            \m_cablesIn[25][14] , \B_int[11] , \m_cablesIn[25][11] , \B_int[12] , 
            \m_cablesIn[25][12] , \B_int[9] , \m_cablesIn[25][9] , \B_int[10] , 
            \m_cablesIn[25][10] , \B_int[7] , \m_cablesIn[25][7] , \B_int[8] , 
            \m_cablesIn[25][8] , \B_int[5] , \m_cablesIn[25][5] , \B_int[6] , 
            \m_cablesIn[25][6] , \B_int[3] , \m_cablesIn[25][3] , \B_int[4] , 
            \m_cablesIn[25][4] , \B_int[1] , \m_cablesIn[25][1] , \B_int[2] , 
            \m_cablesIn[25][2] , \B_int[0] , \frac_div[2] );
    input \m_cablesIn[25][23] ;
    input \QQ_in[25][24] ;
    input GND_net;
    input \m_cablesIn[25][24] ;
    output \QQ_in[26][25] ;
    input \B_int[21] ;
    input \m_cablesIn[25][21] ;
    input \B_int[22] ;
    input \m_cablesIn[25][22] ;
    input \B_int[19] ;
    input \m_cablesIn[25][19] ;
    input \B_int[20] ;
    input \m_cablesIn[25][20] ;
    input \B_int[17] ;
    input \m_cablesIn[25][17] ;
    input \B_int[18] ;
    input \m_cablesIn[25][18] ;
    input \B_int[15] ;
    input \m_cablesIn[25][15] ;
    input \B_int[16] ;
    input \m_cablesIn[25][16] ;
    input \B_int[13] ;
    input \m_cablesIn[25][13] ;
    input \B_int[14] ;
    input \m_cablesIn[25][14] ;
    input \B_int[11] ;
    input \m_cablesIn[25][11] ;
    input \B_int[12] ;
    input \m_cablesIn[25][12] ;
    input \B_int[9] ;
    input \m_cablesIn[25][9] ;
    input \B_int[10] ;
    input \m_cablesIn[25][10] ;
    input \B_int[7] ;
    input \m_cablesIn[25][7] ;
    input \B_int[8] ;
    input \m_cablesIn[25][8] ;
    input \B_int[5] ;
    input \m_cablesIn[25][5] ;
    input \B_int[6] ;
    input \m_cablesIn[25][6] ;
    input \B_int[3] ;
    input \m_cablesIn[25][3] ;
    input \B_int[4] ;
    input \m_cablesIn[25][4] ;
    input \B_int[1] ;
    input \m_cablesIn[25][1] ;
    input \B_int[2] ;
    input \m_cablesIn[25][2] ;
    input \B_int[0] ;
    input \frac_div[2] ;
    
    
    wire n61677, n61676, n61675, n61674, n61673, n61672, n61671, 
        n61670, n61669, n61668, n61667, n61666;
    
    CCU2D add_3745_25 (.A0(\m_cablesIn[25][23] ), .B0(\QQ_in[25][24] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[25][24] ), .B1(\QQ_in[25][24] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n61677), .S1(\QQ_in[26][25] ));
    defparam add_3745_25.INIT0 = 16'h5666;
    defparam add_3745_25.INIT1 = 16'h5999;
    defparam add_3745_25.INJECT1_0 = "NO";
    defparam add_3745_25.INJECT1_1 = "NO";
    CCU2D add_3745_23 (.A0(\B_int[21] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][22] ), 
          .D1(GND_net), .CIN(n61676), .COUT(n61677));
    defparam add_3745_23.INIT0 = 16'h6969;
    defparam add_3745_23.INIT1 = 16'h6969;
    defparam add_3745_23.INJECT1_0 = "NO";
    defparam add_3745_23.INJECT1_1 = "NO";
    CCU2D add_3745_21 (.A0(\B_int[19] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][20] ), 
          .D1(GND_net), .CIN(n61675), .COUT(n61676));
    defparam add_3745_21.INIT0 = 16'h6969;
    defparam add_3745_21.INIT1 = 16'h6969;
    defparam add_3745_21.INJECT1_0 = "NO";
    defparam add_3745_21.INJECT1_1 = "NO";
    CCU2D add_3745_19 (.A0(\B_int[17] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][18] ), 
          .D1(GND_net), .CIN(n61674), .COUT(n61675));
    defparam add_3745_19.INIT0 = 16'h6969;
    defparam add_3745_19.INIT1 = 16'h6969;
    defparam add_3745_19.INJECT1_0 = "NO";
    defparam add_3745_19.INJECT1_1 = "NO";
    CCU2D add_3745_17 (.A0(\B_int[15] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][16] ), 
          .D1(GND_net), .CIN(n61673), .COUT(n61674));
    defparam add_3745_17.INIT0 = 16'h6969;
    defparam add_3745_17.INIT1 = 16'h6969;
    defparam add_3745_17.INJECT1_0 = "NO";
    defparam add_3745_17.INJECT1_1 = "NO";
    CCU2D add_3745_15 (.A0(\B_int[13] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][14] ), 
          .D1(GND_net), .CIN(n61672), .COUT(n61673));
    defparam add_3745_15.INIT0 = 16'h6969;
    defparam add_3745_15.INIT1 = 16'h6969;
    defparam add_3745_15.INJECT1_0 = "NO";
    defparam add_3745_15.INJECT1_1 = "NO";
    CCU2D add_3745_13 (.A0(\B_int[11] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][12] ), 
          .D1(GND_net), .CIN(n61671), .COUT(n61672));
    defparam add_3745_13.INIT0 = 16'h6969;
    defparam add_3745_13.INIT1 = 16'h6969;
    defparam add_3745_13.INJECT1_0 = "NO";
    defparam add_3745_13.INJECT1_1 = "NO";
    CCU2D add_3745_11 (.A0(\B_int[9] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][10] ), 
          .D1(GND_net), .CIN(n61670), .COUT(n61671));
    defparam add_3745_11.INIT0 = 16'h6969;
    defparam add_3745_11.INIT1 = 16'h6969;
    defparam add_3745_11.INJECT1_0 = "NO";
    defparam add_3745_11.INJECT1_1 = "NO";
    CCU2D add_3745_9 (.A0(\B_int[7] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][8] ), 
          .D1(GND_net), .CIN(n61669), .COUT(n61670));
    defparam add_3745_9.INIT0 = 16'h6969;
    defparam add_3745_9.INIT1 = 16'h6969;
    defparam add_3745_9.INJECT1_0 = "NO";
    defparam add_3745_9.INJECT1_1 = "NO";
    CCU2D add_3745_7 (.A0(\B_int[5] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][6] ), 
          .D1(GND_net), .CIN(n61668), .COUT(n61669));
    defparam add_3745_7.INIT0 = 16'h6969;
    defparam add_3745_7.INIT1 = 16'h6969;
    defparam add_3745_7.INJECT1_0 = "NO";
    defparam add_3745_7.INJECT1_1 = "NO";
    CCU2D add_3745_5 (.A0(\B_int[3] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][4] ), 
          .D1(GND_net), .CIN(n61667), .COUT(n61668));
    defparam add_3745_5.INIT0 = 16'h6969;
    defparam add_3745_5.INIT1 = 16'h6969;
    defparam add_3745_5.INJECT1_0 = "NO";
    defparam add_3745_5.INJECT1_1 = "NO";
    CCU2D add_3745_3 (.A0(\B_int[1] ), .B0(\QQ_in[25][24] ), .C0(\m_cablesIn[25][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[25][24] ), .C1(\m_cablesIn[25][2] ), 
          .D1(GND_net), .CIN(n61666), .COUT(n61667));
    defparam add_3745_3.INIT0 = 16'h6969;
    defparam add_3745_3.INIT1 = 16'h6969;
    defparam add_3745_3.INJECT1_0 = "NO";
    defparam add_3745_3.INJECT1_1 = "NO";
    CCU2D add_3745_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[25][24] ), .C1(\frac_div[2] ), .D1(GND_net), 
          .COUT(n61666));
    defparam add_3745_1.INIT0 = 16'hF000;
    defparam add_3745_1.INIT1 = 16'h6969;
    defparam add_3745_1.INJECT1_0 = "NO";
    defparam add_3745_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U8 
//

module \a_s(24)_U8  (\QQ_in[25][24] , \frac_div[2] , \m_cablesIn[24][23] , 
            \QQ_in[24][23] , GND_net, \m_cablesIn[24][24] , \m_cablesIn[25][24] , 
            \B_int[21] , \m_cablesIn[24][21] , \B_int[22] , \m_cablesIn[24][22] , 
            \m_cablesIn[25][22] , \m_cablesIn[25][23] , \B_int[19] , \m_cablesIn[24][19] , 
            \B_int[20] , \m_cablesIn[24][20] , \m_cablesIn[25][20] , \m_cablesIn[25][21] , 
            \B_int[17] , \m_cablesIn[24][17] , \B_int[18] , \m_cablesIn[24][18] , 
            \m_cablesIn[25][18] , \m_cablesIn[25][19] , \B_int[15] , \m_cablesIn[24][15] , 
            \B_int[16] , \m_cablesIn[24][16] , \m_cablesIn[25][16] , \m_cablesIn[25][17] , 
            \B_int[13] , \m_cablesIn[24][13] , \B_int[14] , \m_cablesIn[24][14] , 
            \m_cablesIn[25][14] , \m_cablesIn[25][15] , \B_int[11] , \m_cablesIn[24][11] , 
            \B_int[12] , \m_cablesIn[24][12] , \m_cablesIn[25][12] , \m_cablesIn[25][13] , 
            \B_int[9] , \m_cablesIn[24][9] , \B_int[10] , \m_cablesIn[24][10] , 
            \m_cablesIn[25][10] , \m_cablesIn[25][11] , \B_int[7] , \m_cablesIn[24][7] , 
            \B_int[8] , \m_cablesIn[24][8] , \m_cablesIn[25][8] , \m_cablesIn[25][9] , 
            \B_int[5] , \m_cablesIn[24][5] , \B_int[6] , \m_cablesIn[24][6] , 
            \m_cablesIn[25][6] , \m_cablesIn[25][7] , \B_int[3] , \m_cablesIn[24][3] , 
            \B_int[4] , \m_cablesIn[24][4] , \m_cablesIn[25][4] , \m_cablesIn[25][5] , 
            \B_int[1] , \m_cablesIn[24][1] , \B_int[2] , \m_cablesIn[24][2] , 
            \m_cablesIn[25][2] , \m_cablesIn[25][3] , \B_int[0] , \frac_div[3] , 
            \m_cablesIn[25][1] );
    output \QQ_in[25][24] ;
    output \frac_div[2] ;
    input \m_cablesIn[24][23] ;
    input \QQ_in[24][23] ;
    input GND_net;
    input \m_cablesIn[24][24] ;
    output \m_cablesIn[25][24] ;
    input \B_int[21] ;
    input \m_cablesIn[24][21] ;
    input \B_int[22] ;
    input \m_cablesIn[24][22] ;
    output \m_cablesIn[25][22] ;
    output \m_cablesIn[25][23] ;
    input \B_int[19] ;
    input \m_cablesIn[24][19] ;
    input \B_int[20] ;
    input \m_cablesIn[24][20] ;
    output \m_cablesIn[25][20] ;
    output \m_cablesIn[25][21] ;
    input \B_int[17] ;
    input \m_cablesIn[24][17] ;
    input \B_int[18] ;
    input \m_cablesIn[24][18] ;
    output \m_cablesIn[25][18] ;
    output \m_cablesIn[25][19] ;
    input \B_int[15] ;
    input \m_cablesIn[24][15] ;
    input \B_int[16] ;
    input \m_cablesIn[24][16] ;
    output \m_cablesIn[25][16] ;
    output \m_cablesIn[25][17] ;
    input \B_int[13] ;
    input \m_cablesIn[24][13] ;
    input \B_int[14] ;
    input \m_cablesIn[24][14] ;
    output \m_cablesIn[25][14] ;
    output \m_cablesIn[25][15] ;
    input \B_int[11] ;
    input \m_cablesIn[24][11] ;
    input \B_int[12] ;
    input \m_cablesIn[24][12] ;
    output \m_cablesIn[25][12] ;
    output \m_cablesIn[25][13] ;
    input \B_int[9] ;
    input \m_cablesIn[24][9] ;
    input \B_int[10] ;
    input \m_cablesIn[24][10] ;
    output \m_cablesIn[25][10] ;
    output \m_cablesIn[25][11] ;
    input \B_int[7] ;
    input \m_cablesIn[24][7] ;
    input \B_int[8] ;
    input \m_cablesIn[24][8] ;
    output \m_cablesIn[25][8] ;
    output \m_cablesIn[25][9] ;
    input \B_int[5] ;
    input \m_cablesIn[24][5] ;
    input \B_int[6] ;
    input \m_cablesIn[24][6] ;
    output \m_cablesIn[25][6] ;
    output \m_cablesIn[25][7] ;
    input \B_int[3] ;
    input \m_cablesIn[24][3] ;
    input \B_int[4] ;
    input \m_cablesIn[24][4] ;
    output \m_cablesIn[25][4] ;
    output \m_cablesIn[25][5] ;
    input \B_int[1] ;
    input \m_cablesIn[24][1] ;
    input \B_int[2] ;
    input \m_cablesIn[24][2] ;
    output \m_cablesIn[25][2] ;
    output \m_cablesIn[25][3] ;
    input \B_int[0] ;
    input \frac_div[3] ;
    output \m_cablesIn[25][1] ;
    
    
    wire n61690, n61689, n61688, n61687, n61686, n61685, n61684, 
        n61683, n61682, n61681, n61680, n61679;
    
    LUT4 i3941_1_lut (.A(\QQ_in[25][24] ), .Z(\frac_div[2] )) /* synthesis lut_function=(!(A)) */ ;
    defparam i3941_1_lut.init = 16'h5555;
    CCU2D add_3719_25 (.A0(\m_cablesIn[24][23] ), .B0(\QQ_in[24][23] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[24][24] ), .B1(\QQ_in[24][23] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n61690), .S0(\m_cablesIn[25][24] ), 
          .S1(\QQ_in[25][24] ));
    defparam add_3719_25.INIT0 = 16'h5666;
    defparam add_3719_25.INIT1 = 16'h5999;
    defparam add_3719_25.INJECT1_0 = "NO";
    defparam add_3719_25.INJECT1_1 = "NO";
    CCU2D add_3719_23 (.A0(\B_int[21] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][22] ), 
          .D1(GND_net), .CIN(n61689), .COUT(n61690), .S0(\m_cablesIn[25][22] ), 
          .S1(\m_cablesIn[25][23] ));
    defparam add_3719_23.INIT0 = 16'h6969;
    defparam add_3719_23.INIT1 = 16'h6969;
    defparam add_3719_23.INJECT1_0 = "NO";
    defparam add_3719_23.INJECT1_1 = "NO";
    CCU2D add_3719_21 (.A0(\B_int[19] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][20] ), 
          .D1(GND_net), .CIN(n61688), .COUT(n61689), .S0(\m_cablesIn[25][20] ), 
          .S1(\m_cablesIn[25][21] ));
    defparam add_3719_21.INIT0 = 16'h6969;
    defparam add_3719_21.INIT1 = 16'h6969;
    defparam add_3719_21.INJECT1_0 = "NO";
    defparam add_3719_21.INJECT1_1 = "NO";
    CCU2D add_3719_19 (.A0(\B_int[17] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][18] ), 
          .D1(GND_net), .CIN(n61687), .COUT(n61688), .S0(\m_cablesIn[25][18] ), 
          .S1(\m_cablesIn[25][19] ));
    defparam add_3719_19.INIT0 = 16'h6969;
    defparam add_3719_19.INIT1 = 16'h6969;
    defparam add_3719_19.INJECT1_0 = "NO";
    defparam add_3719_19.INJECT1_1 = "NO";
    CCU2D add_3719_17 (.A0(\B_int[15] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][16] ), 
          .D1(GND_net), .CIN(n61686), .COUT(n61687), .S0(\m_cablesIn[25][16] ), 
          .S1(\m_cablesIn[25][17] ));
    defparam add_3719_17.INIT0 = 16'h6969;
    defparam add_3719_17.INIT1 = 16'h6969;
    defparam add_3719_17.INJECT1_0 = "NO";
    defparam add_3719_17.INJECT1_1 = "NO";
    CCU2D add_3719_15 (.A0(\B_int[13] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][14] ), 
          .D1(GND_net), .CIN(n61685), .COUT(n61686), .S0(\m_cablesIn[25][14] ), 
          .S1(\m_cablesIn[25][15] ));
    defparam add_3719_15.INIT0 = 16'h6969;
    defparam add_3719_15.INIT1 = 16'h6969;
    defparam add_3719_15.INJECT1_0 = "NO";
    defparam add_3719_15.INJECT1_1 = "NO";
    CCU2D add_3719_13 (.A0(\B_int[11] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][12] ), 
          .D1(GND_net), .CIN(n61684), .COUT(n61685), .S0(\m_cablesIn[25][12] ), 
          .S1(\m_cablesIn[25][13] ));
    defparam add_3719_13.INIT0 = 16'h6969;
    defparam add_3719_13.INIT1 = 16'h6969;
    defparam add_3719_13.INJECT1_0 = "NO";
    defparam add_3719_13.INJECT1_1 = "NO";
    CCU2D add_3719_11 (.A0(\B_int[9] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][10] ), 
          .D1(GND_net), .CIN(n61683), .COUT(n61684), .S0(\m_cablesIn[25][10] ), 
          .S1(\m_cablesIn[25][11] ));
    defparam add_3719_11.INIT0 = 16'h6969;
    defparam add_3719_11.INIT1 = 16'h6969;
    defparam add_3719_11.INJECT1_0 = "NO";
    defparam add_3719_11.INJECT1_1 = "NO";
    CCU2D add_3719_9 (.A0(\B_int[7] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][8] ), 
          .D1(GND_net), .CIN(n61682), .COUT(n61683), .S0(\m_cablesIn[25][8] ), 
          .S1(\m_cablesIn[25][9] ));
    defparam add_3719_9.INIT0 = 16'h6969;
    defparam add_3719_9.INIT1 = 16'h6969;
    defparam add_3719_9.INJECT1_0 = "NO";
    defparam add_3719_9.INJECT1_1 = "NO";
    CCU2D add_3719_7 (.A0(\B_int[5] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][6] ), 
          .D1(GND_net), .CIN(n61681), .COUT(n61682), .S0(\m_cablesIn[25][6] ), 
          .S1(\m_cablesIn[25][7] ));
    defparam add_3719_7.INIT0 = 16'h6969;
    defparam add_3719_7.INIT1 = 16'h6969;
    defparam add_3719_7.INJECT1_0 = "NO";
    defparam add_3719_7.INJECT1_1 = "NO";
    CCU2D add_3719_5 (.A0(\B_int[3] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][4] ), 
          .D1(GND_net), .CIN(n61680), .COUT(n61681), .S0(\m_cablesIn[25][4] ), 
          .S1(\m_cablesIn[25][5] ));
    defparam add_3719_5.INIT0 = 16'h6969;
    defparam add_3719_5.INIT1 = 16'h6969;
    defparam add_3719_5.INJECT1_0 = "NO";
    defparam add_3719_5.INJECT1_1 = "NO";
    CCU2D add_3719_3 (.A0(\B_int[1] ), .B0(\QQ_in[24][23] ), .C0(\m_cablesIn[24][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[24][23] ), .C1(\m_cablesIn[24][2] ), 
          .D1(GND_net), .CIN(n61679), .COUT(n61680), .S0(\m_cablesIn[25][2] ), 
          .S1(\m_cablesIn[25][3] ));
    defparam add_3719_3.INIT0 = 16'h6969;
    defparam add_3719_3.INIT1 = 16'h6969;
    defparam add_3719_3.INJECT1_0 = "NO";
    defparam add_3719_3.INJECT1_1 = "NO";
    CCU2D add_3719_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[24][23] ), .C1(\frac_div[3] ), .D1(GND_net), 
          .COUT(n61679), .S1(\m_cablesIn[25][1] ));
    defparam add_3719_1.INIT0 = 16'hF000;
    defparam add_3719_1.INIT1 = 16'h6969;
    defparam add_3719_1.INJECT1_0 = "NO";
    defparam add_3719_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U9 
//

module \a_s(24)_U9  (\m_cablesIn[23][23] , \QQ_in[23][22] , GND_net, \m_cablesIn[23][24] , 
            \m_cablesIn[24][24] , \QQ_in[24][23] , \B_int[21] , \m_cablesIn[23][21] , 
            \B_int[22] , \m_cablesIn[23][22] , \m_cablesIn[24][22] , \m_cablesIn[24][23] , 
            \B_int[19] , \m_cablesIn[23][19] , \B_int[20] , \m_cablesIn[23][20] , 
            \m_cablesIn[24][20] , \m_cablesIn[24][21] , \B_int[17] , \m_cablesIn[23][17] , 
            \B_int[18] , \m_cablesIn[23][18] , \m_cablesIn[24][18] , \m_cablesIn[24][19] , 
            \B_int[15] , \m_cablesIn[23][15] , \B_int[16] , \m_cablesIn[23][16] , 
            \m_cablesIn[24][16] , \m_cablesIn[24][17] , \B_int[13] , \m_cablesIn[23][13] , 
            \B_int[14] , \m_cablesIn[23][14] , \m_cablesIn[24][14] , \m_cablesIn[24][15] , 
            \B_int[11] , \m_cablesIn[23][11] , \B_int[12] , \m_cablesIn[23][12] , 
            \m_cablesIn[24][12] , \m_cablesIn[24][13] , \B_int[9] , \m_cablesIn[23][9] , 
            \B_int[10] , \m_cablesIn[23][10] , \m_cablesIn[24][10] , \m_cablesIn[24][11] , 
            \B_int[7] , \m_cablesIn[23][7] , \B_int[8] , \m_cablesIn[23][8] , 
            \m_cablesIn[24][8] , \m_cablesIn[24][9] , \B_int[5] , \m_cablesIn[23][5] , 
            \B_int[6] , \m_cablesIn[23][6] , \m_cablesIn[24][6] , \m_cablesIn[24][7] , 
            \B_int[3] , \m_cablesIn[23][3] , \B_int[4] , \m_cablesIn[23][4] , 
            \m_cablesIn[24][4] , \m_cablesIn[24][5] , \B_int[1] , \m_cablesIn[23][1] , 
            \B_int[2] , \m_cablesIn[23][2] , \m_cablesIn[24][2] , \m_cablesIn[24][3] , 
            \B_int[0] , \frac_div[4] , \m_cablesIn[24][1] );
    input \m_cablesIn[23][23] ;
    input \QQ_in[23][22] ;
    input GND_net;
    input \m_cablesIn[23][24] ;
    output \m_cablesIn[24][24] ;
    output \QQ_in[24][23] ;
    input \B_int[21] ;
    input \m_cablesIn[23][21] ;
    input \B_int[22] ;
    input \m_cablesIn[23][22] ;
    output \m_cablesIn[24][22] ;
    output \m_cablesIn[24][23] ;
    input \B_int[19] ;
    input \m_cablesIn[23][19] ;
    input \B_int[20] ;
    input \m_cablesIn[23][20] ;
    output \m_cablesIn[24][20] ;
    output \m_cablesIn[24][21] ;
    input \B_int[17] ;
    input \m_cablesIn[23][17] ;
    input \B_int[18] ;
    input \m_cablesIn[23][18] ;
    output \m_cablesIn[24][18] ;
    output \m_cablesIn[24][19] ;
    input \B_int[15] ;
    input \m_cablesIn[23][15] ;
    input \B_int[16] ;
    input \m_cablesIn[23][16] ;
    output \m_cablesIn[24][16] ;
    output \m_cablesIn[24][17] ;
    input \B_int[13] ;
    input \m_cablesIn[23][13] ;
    input \B_int[14] ;
    input \m_cablesIn[23][14] ;
    output \m_cablesIn[24][14] ;
    output \m_cablesIn[24][15] ;
    input \B_int[11] ;
    input \m_cablesIn[23][11] ;
    input \B_int[12] ;
    input \m_cablesIn[23][12] ;
    output \m_cablesIn[24][12] ;
    output \m_cablesIn[24][13] ;
    input \B_int[9] ;
    input \m_cablesIn[23][9] ;
    input \B_int[10] ;
    input \m_cablesIn[23][10] ;
    output \m_cablesIn[24][10] ;
    output \m_cablesIn[24][11] ;
    input \B_int[7] ;
    input \m_cablesIn[23][7] ;
    input \B_int[8] ;
    input \m_cablesIn[23][8] ;
    output \m_cablesIn[24][8] ;
    output \m_cablesIn[24][9] ;
    input \B_int[5] ;
    input \m_cablesIn[23][5] ;
    input \B_int[6] ;
    input \m_cablesIn[23][6] ;
    output \m_cablesIn[24][6] ;
    output \m_cablesIn[24][7] ;
    input \B_int[3] ;
    input \m_cablesIn[23][3] ;
    input \B_int[4] ;
    input \m_cablesIn[23][4] ;
    output \m_cablesIn[24][4] ;
    output \m_cablesIn[24][5] ;
    input \B_int[1] ;
    input \m_cablesIn[23][1] ;
    input \B_int[2] ;
    input \m_cablesIn[23][2] ;
    output \m_cablesIn[24][2] ;
    output \m_cablesIn[24][3] ;
    input \B_int[0] ;
    input \frac_div[4] ;
    output \m_cablesIn[24][1] ;
    
    
    wire n62230, n62229, n62228, n62227, n62226, n62225, n62224, 
        n62223, n62222, n62221, n62220, n62219;
    
    CCU2D add_3693_25 (.A0(\m_cablesIn[23][23] ), .B0(\QQ_in[23][22] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[23][24] ), .B1(\QQ_in[23][22] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62230), .S0(\m_cablesIn[24][24] ), 
          .S1(\QQ_in[24][23] ));
    defparam add_3693_25.INIT0 = 16'h5666;
    defparam add_3693_25.INIT1 = 16'h5999;
    defparam add_3693_25.INJECT1_0 = "NO";
    defparam add_3693_25.INJECT1_1 = "NO";
    CCU2D add_3693_23 (.A0(\B_int[21] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][22] ), 
          .D1(GND_net), .CIN(n62229), .COUT(n62230), .S0(\m_cablesIn[24][22] ), 
          .S1(\m_cablesIn[24][23] ));
    defparam add_3693_23.INIT0 = 16'h6969;
    defparam add_3693_23.INIT1 = 16'h6969;
    defparam add_3693_23.INJECT1_0 = "NO";
    defparam add_3693_23.INJECT1_1 = "NO";
    CCU2D add_3693_21 (.A0(\B_int[19] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][20] ), 
          .D1(GND_net), .CIN(n62228), .COUT(n62229), .S0(\m_cablesIn[24][20] ), 
          .S1(\m_cablesIn[24][21] ));
    defparam add_3693_21.INIT0 = 16'h6969;
    defparam add_3693_21.INIT1 = 16'h6969;
    defparam add_3693_21.INJECT1_0 = "NO";
    defparam add_3693_21.INJECT1_1 = "NO";
    CCU2D add_3693_19 (.A0(\B_int[17] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][18] ), 
          .D1(GND_net), .CIN(n62227), .COUT(n62228), .S0(\m_cablesIn[24][18] ), 
          .S1(\m_cablesIn[24][19] ));
    defparam add_3693_19.INIT0 = 16'h6969;
    defparam add_3693_19.INIT1 = 16'h6969;
    defparam add_3693_19.INJECT1_0 = "NO";
    defparam add_3693_19.INJECT1_1 = "NO";
    CCU2D add_3693_17 (.A0(\B_int[15] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][16] ), 
          .D1(GND_net), .CIN(n62226), .COUT(n62227), .S0(\m_cablesIn[24][16] ), 
          .S1(\m_cablesIn[24][17] ));
    defparam add_3693_17.INIT0 = 16'h6969;
    defparam add_3693_17.INIT1 = 16'h6969;
    defparam add_3693_17.INJECT1_0 = "NO";
    defparam add_3693_17.INJECT1_1 = "NO";
    CCU2D add_3693_15 (.A0(\B_int[13] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][14] ), 
          .D1(GND_net), .CIN(n62225), .COUT(n62226), .S0(\m_cablesIn[24][14] ), 
          .S1(\m_cablesIn[24][15] ));
    defparam add_3693_15.INIT0 = 16'h6969;
    defparam add_3693_15.INIT1 = 16'h6969;
    defparam add_3693_15.INJECT1_0 = "NO";
    defparam add_3693_15.INJECT1_1 = "NO";
    CCU2D add_3693_13 (.A0(\B_int[11] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][12] ), 
          .D1(GND_net), .CIN(n62224), .COUT(n62225), .S0(\m_cablesIn[24][12] ), 
          .S1(\m_cablesIn[24][13] ));
    defparam add_3693_13.INIT0 = 16'h6969;
    defparam add_3693_13.INIT1 = 16'h6969;
    defparam add_3693_13.INJECT1_0 = "NO";
    defparam add_3693_13.INJECT1_1 = "NO";
    CCU2D add_3693_11 (.A0(\B_int[9] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][10] ), 
          .D1(GND_net), .CIN(n62223), .COUT(n62224), .S0(\m_cablesIn[24][10] ), 
          .S1(\m_cablesIn[24][11] ));
    defparam add_3693_11.INIT0 = 16'h6969;
    defparam add_3693_11.INIT1 = 16'h6969;
    defparam add_3693_11.INJECT1_0 = "NO";
    defparam add_3693_11.INJECT1_1 = "NO";
    CCU2D add_3693_9 (.A0(\B_int[7] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][8] ), 
          .D1(GND_net), .CIN(n62222), .COUT(n62223), .S0(\m_cablesIn[24][8] ), 
          .S1(\m_cablesIn[24][9] ));
    defparam add_3693_9.INIT0 = 16'h6969;
    defparam add_3693_9.INIT1 = 16'h6969;
    defparam add_3693_9.INJECT1_0 = "NO";
    defparam add_3693_9.INJECT1_1 = "NO";
    CCU2D add_3693_7 (.A0(\B_int[5] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][6] ), 
          .D1(GND_net), .CIN(n62221), .COUT(n62222), .S0(\m_cablesIn[24][6] ), 
          .S1(\m_cablesIn[24][7] ));
    defparam add_3693_7.INIT0 = 16'h6969;
    defparam add_3693_7.INIT1 = 16'h6969;
    defparam add_3693_7.INJECT1_0 = "NO";
    defparam add_3693_7.INJECT1_1 = "NO";
    CCU2D add_3693_5 (.A0(\B_int[3] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][4] ), 
          .D1(GND_net), .CIN(n62220), .COUT(n62221), .S0(\m_cablesIn[24][4] ), 
          .S1(\m_cablesIn[24][5] ));
    defparam add_3693_5.INIT0 = 16'h6969;
    defparam add_3693_5.INIT1 = 16'h6969;
    defparam add_3693_5.INJECT1_0 = "NO";
    defparam add_3693_5.INJECT1_1 = "NO";
    CCU2D add_3693_3 (.A0(\B_int[1] ), .B0(\QQ_in[23][22] ), .C0(\m_cablesIn[23][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[23][22] ), .C1(\m_cablesIn[23][2] ), 
          .D1(GND_net), .CIN(n62219), .COUT(n62220), .S0(\m_cablesIn[24][2] ), 
          .S1(\m_cablesIn[24][3] ));
    defparam add_3693_3.INIT0 = 16'h6969;
    defparam add_3693_3.INIT1 = 16'h6969;
    defparam add_3693_3.INJECT1_0 = "NO";
    defparam add_3693_3.INJECT1_1 = "NO";
    CCU2D add_3693_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[23][22] ), .C1(\frac_div[4] ), .D1(GND_net), 
          .COUT(n62219), .S1(\m_cablesIn[24][1] ));
    defparam add_3693_1.INIT0 = 16'hF000;
    defparam add_3693_1.INIT1 = 16'h6969;
    defparam add_3693_1.INJECT1_0 = "NO";
    defparam add_3693_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U10 
//

module \a_s(24)_U10  (\m_cablesIn[22][23] , \QQ_in[22][21] , GND_net, 
            \m_cablesIn[22][24] , \m_cablesIn[23][24] , \QQ_in[23][22] , 
            \B_int[21] , \m_cablesIn[22][21] , \B_int[22] , \m_cablesIn[22][22] , 
            \m_cablesIn[23][22] , \m_cablesIn[23][23] , \B_int[19] , \m_cablesIn[22][19] , 
            \B_int[20] , \m_cablesIn[22][20] , \m_cablesIn[23][20] , \m_cablesIn[23][21] , 
            \B_int[17] , \m_cablesIn[22][17] , \B_int[18] , \m_cablesIn[22][18] , 
            \m_cablesIn[23][18] , \m_cablesIn[23][19] , \B_int[15] , \m_cablesIn[22][15] , 
            \B_int[16] , \m_cablesIn[22][16] , \m_cablesIn[23][16] , \m_cablesIn[23][17] , 
            \B_int[13] , \m_cablesIn[22][13] , \B_int[14] , \m_cablesIn[22][14] , 
            \m_cablesIn[23][14] , \m_cablesIn[23][15] , \B_int[11] , \m_cablesIn[22][11] , 
            \B_int[12] , \m_cablesIn[22][12] , \m_cablesIn[23][12] , \m_cablesIn[23][13] , 
            \B_int[9] , \m_cablesIn[22][9] , \B_int[10] , \m_cablesIn[22][10] , 
            \m_cablesIn[23][10] , \m_cablesIn[23][11] , \B_int[7] , \m_cablesIn[22][7] , 
            \B_int[8] , \m_cablesIn[22][8] , \m_cablesIn[23][8] , \m_cablesIn[23][9] , 
            \B_int[5] , \m_cablesIn[22][5] , \B_int[6] , \m_cablesIn[22][6] , 
            \m_cablesIn[23][6] , \m_cablesIn[23][7] , \B_int[3] , \m_cablesIn[22][3] , 
            \B_int[4] , \m_cablesIn[22][4] , \m_cablesIn[23][4] , \m_cablesIn[23][5] , 
            \B_int[1] , \m_cablesIn[22][1] , \B_int[2] , \m_cablesIn[22][2] , 
            \m_cablesIn[23][2] , \m_cablesIn[23][3] , \B_int[0] , \frac_div[5] , 
            \m_cablesIn[23][1] );
    input \m_cablesIn[22][23] ;
    input \QQ_in[22][21] ;
    input GND_net;
    input \m_cablesIn[22][24] ;
    output \m_cablesIn[23][24] ;
    output \QQ_in[23][22] ;
    input \B_int[21] ;
    input \m_cablesIn[22][21] ;
    input \B_int[22] ;
    input \m_cablesIn[22][22] ;
    output \m_cablesIn[23][22] ;
    output \m_cablesIn[23][23] ;
    input \B_int[19] ;
    input \m_cablesIn[22][19] ;
    input \B_int[20] ;
    input \m_cablesIn[22][20] ;
    output \m_cablesIn[23][20] ;
    output \m_cablesIn[23][21] ;
    input \B_int[17] ;
    input \m_cablesIn[22][17] ;
    input \B_int[18] ;
    input \m_cablesIn[22][18] ;
    output \m_cablesIn[23][18] ;
    output \m_cablesIn[23][19] ;
    input \B_int[15] ;
    input \m_cablesIn[22][15] ;
    input \B_int[16] ;
    input \m_cablesIn[22][16] ;
    output \m_cablesIn[23][16] ;
    output \m_cablesIn[23][17] ;
    input \B_int[13] ;
    input \m_cablesIn[22][13] ;
    input \B_int[14] ;
    input \m_cablesIn[22][14] ;
    output \m_cablesIn[23][14] ;
    output \m_cablesIn[23][15] ;
    input \B_int[11] ;
    input \m_cablesIn[22][11] ;
    input \B_int[12] ;
    input \m_cablesIn[22][12] ;
    output \m_cablesIn[23][12] ;
    output \m_cablesIn[23][13] ;
    input \B_int[9] ;
    input \m_cablesIn[22][9] ;
    input \B_int[10] ;
    input \m_cablesIn[22][10] ;
    output \m_cablesIn[23][10] ;
    output \m_cablesIn[23][11] ;
    input \B_int[7] ;
    input \m_cablesIn[22][7] ;
    input \B_int[8] ;
    input \m_cablesIn[22][8] ;
    output \m_cablesIn[23][8] ;
    output \m_cablesIn[23][9] ;
    input \B_int[5] ;
    input \m_cablesIn[22][5] ;
    input \B_int[6] ;
    input \m_cablesIn[22][6] ;
    output \m_cablesIn[23][6] ;
    output \m_cablesIn[23][7] ;
    input \B_int[3] ;
    input \m_cablesIn[22][3] ;
    input \B_int[4] ;
    input \m_cablesIn[22][4] ;
    output \m_cablesIn[23][4] ;
    output \m_cablesIn[23][5] ;
    input \B_int[1] ;
    input \m_cablesIn[22][1] ;
    input \B_int[2] ;
    input \m_cablesIn[22][2] ;
    output \m_cablesIn[23][2] ;
    output \m_cablesIn[23][3] ;
    input \B_int[0] ;
    input \frac_div[5] ;
    output \m_cablesIn[23][1] ;
    
    
    wire n62243, n62242, n62241, n62240, n62239, n62238, n62237, 
        n62236, n62235, n62234, n62233, n62232;
    
    CCU2D add_3667_25 (.A0(\m_cablesIn[22][23] ), .B0(\QQ_in[22][21] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[22][24] ), .B1(\QQ_in[22][21] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62243), .S0(\m_cablesIn[23][24] ), 
          .S1(\QQ_in[23][22] ));
    defparam add_3667_25.INIT0 = 16'h5666;
    defparam add_3667_25.INIT1 = 16'h5999;
    defparam add_3667_25.INJECT1_0 = "NO";
    defparam add_3667_25.INJECT1_1 = "NO";
    CCU2D add_3667_23 (.A0(\B_int[21] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][22] ), 
          .D1(GND_net), .CIN(n62242), .COUT(n62243), .S0(\m_cablesIn[23][22] ), 
          .S1(\m_cablesIn[23][23] ));
    defparam add_3667_23.INIT0 = 16'h6969;
    defparam add_3667_23.INIT1 = 16'h6969;
    defparam add_3667_23.INJECT1_0 = "NO";
    defparam add_3667_23.INJECT1_1 = "NO";
    CCU2D add_3667_21 (.A0(\B_int[19] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][20] ), 
          .D1(GND_net), .CIN(n62241), .COUT(n62242), .S0(\m_cablesIn[23][20] ), 
          .S1(\m_cablesIn[23][21] ));
    defparam add_3667_21.INIT0 = 16'h6969;
    defparam add_3667_21.INIT1 = 16'h6969;
    defparam add_3667_21.INJECT1_0 = "NO";
    defparam add_3667_21.INJECT1_1 = "NO";
    CCU2D add_3667_19 (.A0(\B_int[17] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][18] ), 
          .D1(GND_net), .CIN(n62240), .COUT(n62241), .S0(\m_cablesIn[23][18] ), 
          .S1(\m_cablesIn[23][19] ));
    defparam add_3667_19.INIT0 = 16'h6969;
    defparam add_3667_19.INIT1 = 16'h6969;
    defparam add_3667_19.INJECT1_0 = "NO";
    defparam add_3667_19.INJECT1_1 = "NO";
    CCU2D add_3667_17 (.A0(\B_int[15] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][16] ), 
          .D1(GND_net), .CIN(n62239), .COUT(n62240), .S0(\m_cablesIn[23][16] ), 
          .S1(\m_cablesIn[23][17] ));
    defparam add_3667_17.INIT0 = 16'h6969;
    defparam add_3667_17.INIT1 = 16'h6969;
    defparam add_3667_17.INJECT1_0 = "NO";
    defparam add_3667_17.INJECT1_1 = "NO";
    CCU2D add_3667_15 (.A0(\B_int[13] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][14] ), 
          .D1(GND_net), .CIN(n62238), .COUT(n62239), .S0(\m_cablesIn[23][14] ), 
          .S1(\m_cablesIn[23][15] ));
    defparam add_3667_15.INIT0 = 16'h6969;
    defparam add_3667_15.INIT1 = 16'h6969;
    defparam add_3667_15.INJECT1_0 = "NO";
    defparam add_3667_15.INJECT1_1 = "NO";
    CCU2D add_3667_13 (.A0(\B_int[11] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][12] ), 
          .D1(GND_net), .CIN(n62237), .COUT(n62238), .S0(\m_cablesIn[23][12] ), 
          .S1(\m_cablesIn[23][13] ));
    defparam add_3667_13.INIT0 = 16'h6969;
    defparam add_3667_13.INIT1 = 16'h6969;
    defparam add_3667_13.INJECT1_0 = "NO";
    defparam add_3667_13.INJECT1_1 = "NO";
    CCU2D add_3667_11 (.A0(\B_int[9] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][10] ), 
          .D1(GND_net), .CIN(n62236), .COUT(n62237), .S0(\m_cablesIn[23][10] ), 
          .S1(\m_cablesIn[23][11] ));
    defparam add_3667_11.INIT0 = 16'h6969;
    defparam add_3667_11.INIT1 = 16'h6969;
    defparam add_3667_11.INJECT1_0 = "NO";
    defparam add_3667_11.INJECT1_1 = "NO";
    CCU2D add_3667_9 (.A0(\B_int[7] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][8] ), 
          .D1(GND_net), .CIN(n62235), .COUT(n62236), .S0(\m_cablesIn[23][8] ), 
          .S1(\m_cablesIn[23][9] ));
    defparam add_3667_9.INIT0 = 16'h6969;
    defparam add_3667_9.INIT1 = 16'h6969;
    defparam add_3667_9.INJECT1_0 = "NO";
    defparam add_3667_9.INJECT1_1 = "NO";
    CCU2D add_3667_7 (.A0(\B_int[5] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][6] ), 
          .D1(GND_net), .CIN(n62234), .COUT(n62235), .S0(\m_cablesIn[23][6] ), 
          .S1(\m_cablesIn[23][7] ));
    defparam add_3667_7.INIT0 = 16'h6969;
    defparam add_3667_7.INIT1 = 16'h6969;
    defparam add_3667_7.INJECT1_0 = "NO";
    defparam add_3667_7.INJECT1_1 = "NO";
    CCU2D add_3667_5 (.A0(\B_int[3] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][4] ), 
          .D1(GND_net), .CIN(n62233), .COUT(n62234), .S0(\m_cablesIn[23][4] ), 
          .S1(\m_cablesIn[23][5] ));
    defparam add_3667_5.INIT0 = 16'h6969;
    defparam add_3667_5.INIT1 = 16'h6969;
    defparam add_3667_5.INJECT1_0 = "NO";
    defparam add_3667_5.INJECT1_1 = "NO";
    CCU2D add_3667_3 (.A0(\B_int[1] ), .B0(\QQ_in[22][21] ), .C0(\m_cablesIn[22][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[22][21] ), .C1(\m_cablesIn[22][2] ), 
          .D1(GND_net), .CIN(n62232), .COUT(n62233), .S0(\m_cablesIn[23][2] ), 
          .S1(\m_cablesIn[23][3] ));
    defparam add_3667_3.INIT0 = 16'h6969;
    defparam add_3667_3.INIT1 = 16'h6969;
    defparam add_3667_3.INJECT1_0 = "NO";
    defparam add_3667_3.INJECT1_1 = "NO";
    CCU2D add_3667_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[22][21] ), .C1(\frac_div[5] ), .D1(GND_net), 
          .COUT(n62232), .S1(\m_cablesIn[23][1] ));
    defparam add_3667_1.INIT0 = 16'hF000;
    defparam add_3667_1.INIT1 = 16'h6969;
    defparam add_3667_1.INJECT1_0 = "NO";
    defparam add_3667_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U11 
//

module \a_s(24)_U11  (\m_cablesIn[21][23] , \QQ_in[21][20] , GND_net, 
            \m_cablesIn[21][24] , \m_cablesIn[22][24] , \QQ_in[22][21] , 
            \B_int[21] , \m_cablesIn[21][21] , \B_int[22] , \m_cablesIn[21][22] , 
            \m_cablesIn[22][22] , \m_cablesIn[22][23] , \B_int[19] , \m_cablesIn[21][19] , 
            \B_int[20] , \m_cablesIn[21][20] , \m_cablesIn[22][20] , \m_cablesIn[22][21] , 
            \B_int[17] , \m_cablesIn[21][17] , \B_int[18] , \m_cablesIn[21][18] , 
            \m_cablesIn[22][18] , \m_cablesIn[22][19] , \B_int[15] , \m_cablesIn[21][15] , 
            \B_int[16] , \m_cablesIn[21][16] , \m_cablesIn[22][16] , \m_cablesIn[22][17] , 
            \B_int[13] , \m_cablesIn[21][13] , \B_int[14] , \m_cablesIn[21][14] , 
            \m_cablesIn[22][14] , \m_cablesIn[22][15] , \B_int[11] , \m_cablesIn[21][11] , 
            \B_int[12] , \m_cablesIn[21][12] , \m_cablesIn[22][12] , \m_cablesIn[22][13] , 
            \B_int[9] , \m_cablesIn[21][9] , \B_int[10] , \m_cablesIn[21][10] , 
            \m_cablesIn[22][10] , \m_cablesIn[22][11] , \B_int[7] , \m_cablesIn[21][7] , 
            \B_int[8] , \m_cablesIn[21][8] , \m_cablesIn[22][8] , \m_cablesIn[22][9] , 
            \B_int[5] , \m_cablesIn[21][5] , \B_int[6] , \m_cablesIn[21][6] , 
            \m_cablesIn[22][6] , \m_cablesIn[22][7] , \B_int[3] , \m_cablesIn[21][3] , 
            \B_int[4] , \m_cablesIn[21][4] , \m_cablesIn[22][4] , \m_cablesIn[22][5] , 
            \B_int[1] , \m_cablesIn[21][1] , \B_int[2] , \m_cablesIn[21][2] , 
            \m_cablesIn[22][2] , \m_cablesIn[22][3] , \B_int[0] , \frac_div[6] , 
            \m_cablesIn[22][1] );
    input \m_cablesIn[21][23] ;
    input \QQ_in[21][20] ;
    input GND_net;
    input \m_cablesIn[21][24] ;
    output \m_cablesIn[22][24] ;
    output \QQ_in[22][21] ;
    input \B_int[21] ;
    input \m_cablesIn[21][21] ;
    input \B_int[22] ;
    input \m_cablesIn[21][22] ;
    output \m_cablesIn[22][22] ;
    output \m_cablesIn[22][23] ;
    input \B_int[19] ;
    input \m_cablesIn[21][19] ;
    input \B_int[20] ;
    input \m_cablesIn[21][20] ;
    output \m_cablesIn[22][20] ;
    output \m_cablesIn[22][21] ;
    input \B_int[17] ;
    input \m_cablesIn[21][17] ;
    input \B_int[18] ;
    input \m_cablesIn[21][18] ;
    output \m_cablesIn[22][18] ;
    output \m_cablesIn[22][19] ;
    input \B_int[15] ;
    input \m_cablesIn[21][15] ;
    input \B_int[16] ;
    input \m_cablesIn[21][16] ;
    output \m_cablesIn[22][16] ;
    output \m_cablesIn[22][17] ;
    input \B_int[13] ;
    input \m_cablesIn[21][13] ;
    input \B_int[14] ;
    input \m_cablesIn[21][14] ;
    output \m_cablesIn[22][14] ;
    output \m_cablesIn[22][15] ;
    input \B_int[11] ;
    input \m_cablesIn[21][11] ;
    input \B_int[12] ;
    input \m_cablesIn[21][12] ;
    output \m_cablesIn[22][12] ;
    output \m_cablesIn[22][13] ;
    input \B_int[9] ;
    input \m_cablesIn[21][9] ;
    input \B_int[10] ;
    input \m_cablesIn[21][10] ;
    output \m_cablesIn[22][10] ;
    output \m_cablesIn[22][11] ;
    input \B_int[7] ;
    input \m_cablesIn[21][7] ;
    input \B_int[8] ;
    input \m_cablesIn[21][8] ;
    output \m_cablesIn[22][8] ;
    output \m_cablesIn[22][9] ;
    input \B_int[5] ;
    input \m_cablesIn[21][5] ;
    input \B_int[6] ;
    input \m_cablesIn[21][6] ;
    output \m_cablesIn[22][6] ;
    output \m_cablesIn[22][7] ;
    input \B_int[3] ;
    input \m_cablesIn[21][3] ;
    input \B_int[4] ;
    input \m_cablesIn[21][4] ;
    output \m_cablesIn[22][4] ;
    output \m_cablesIn[22][5] ;
    input \B_int[1] ;
    input \m_cablesIn[21][1] ;
    input \B_int[2] ;
    input \m_cablesIn[21][2] ;
    output \m_cablesIn[22][2] ;
    output \m_cablesIn[22][3] ;
    input \B_int[0] ;
    input \frac_div[6] ;
    output \m_cablesIn[22][1] ;
    
    
    wire n62256, n62255, n62254, n62253, n62252, n62251, n62250, 
        n62249, n62248, n62247, n62246, n62245;
    
    CCU2D add_3641_25 (.A0(\m_cablesIn[21][23] ), .B0(\QQ_in[21][20] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[21][24] ), .B1(\QQ_in[21][20] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62256), .S0(\m_cablesIn[22][24] ), 
          .S1(\QQ_in[22][21] ));
    defparam add_3641_25.INIT0 = 16'h5666;
    defparam add_3641_25.INIT1 = 16'h5999;
    defparam add_3641_25.INJECT1_0 = "NO";
    defparam add_3641_25.INJECT1_1 = "NO";
    CCU2D add_3641_23 (.A0(\B_int[21] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][22] ), 
          .D1(GND_net), .CIN(n62255), .COUT(n62256), .S0(\m_cablesIn[22][22] ), 
          .S1(\m_cablesIn[22][23] ));
    defparam add_3641_23.INIT0 = 16'h6969;
    defparam add_3641_23.INIT1 = 16'h6969;
    defparam add_3641_23.INJECT1_0 = "NO";
    defparam add_3641_23.INJECT1_1 = "NO";
    CCU2D add_3641_21 (.A0(\B_int[19] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][20] ), 
          .D1(GND_net), .CIN(n62254), .COUT(n62255), .S0(\m_cablesIn[22][20] ), 
          .S1(\m_cablesIn[22][21] ));
    defparam add_3641_21.INIT0 = 16'h6969;
    defparam add_3641_21.INIT1 = 16'h6969;
    defparam add_3641_21.INJECT1_0 = "NO";
    defparam add_3641_21.INJECT1_1 = "NO";
    CCU2D add_3641_19 (.A0(\B_int[17] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][18] ), 
          .D1(GND_net), .CIN(n62253), .COUT(n62254), .S0(\m_cablesIn[22][18] ), 
          .S1(\m_cablesIn[22][19] ));
    defparam add_3641_19.INIT0 = 16'h6969;
    defparam add_3641_19.INIT1 = 16'h6969;
    defparam add_3641_19.INJECT1_0 = "NO";
    defparam add_3641_19.INJECT1_1 = "NO";
    CCU2D add_3641_17 (.A0(\B_int[15] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][16] ), 
          .D1(GND_net), .CIN(n62252), .COUT(n62253), .S0(\m_cablesIn[22][16] ), 
          .S1(\m_cablesIn[22][17] ));
    defparam add_3641_17.INIT0 = 16'h6969;
    defparam add_3641_17.INIT1 = 16'h6969;
    defparam add_3641_17.INJECT1_0 = "NO";
    defparam add_3641_17.INJECT1_1 = "NO";
    CCU2D add_3641_15 (.A0(\B_int[13] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][14] ), 
          .D1(GND_net), .CIN(n62251), .COUT(n62252), .S0(\m_cablesIn[22][14] ), 
          .S1(\m_cablesIn[22][15] ));
    defparam add_3641_15.INIT0 = 16'h6969;
    defparam add_3641_15.INIT1 = 16'h6969;
    defparam add_3641_15.INJECT1_0 = "NO";
    defparam add_3641_15.INJECT1_1 = "NO";
    CCU2D add_3641_13 (.A0(\B_int[11] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][12] ), 
          .D1(GND_net), .CIN(n62250), .COUT(n62251), .S0(\m_cablesIn[22][12] ), 
          .S1(\m_cablesIn[22][13] ));
    defparam add_3641_13.INIT0 = 16'h6969;
    defparam add_3641_13.INIT1 = 16'h6969;
    defparam add_3641_13.INJECT1_0 = "NO";
    defparam add_3641_13.INJECT1_1 = "NO";
    CCU2D add_3641_11 (.A0(\B_int[9] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][10] ), 
          .D1(GND_net), .CIN(n62249), .COUT(n62250), .S0(\m_cablesIn[22][10] ), 
          .S1(\m_cablesIn[22][11] ));
    defparam add_3641_11.INIT0 = 16'h6969;
    defparam add_3641_11.INIT1 = 16'h6969;
    defparam add_3641_11.INJECT1_0 = "NO";
    defparam add_3641_11.INJECT1_1 = "NO";
    CCU2D add_3641_9 (.A0(\B_int[7] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][8] ), 
          .D1(GND_net), .CIN(n62248), .COUT(n62249), .S0(\m_cablesIn[22][8] ), 
          .S1(\m_cablesIn[22][9] ));
    defparam add_3641_9.INIT0 = 16'h6969;
    defparam add_3641_9.INIT1 = 16'h6969;
    defparam add_3641_9.INJECT1_0 = "NO";
    defparam add_3641_9.INJECT1_1 = "NO";
    CCU2D add_3641_7 (.A0(\B_int[5] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][6] ), 
          .D1(GND_net), .CIN(n62247), .COUT(n62248), .S0(\m_cablesIn[22][6] ), 
          .S1(\m_cablesIn[22][7] ));
    defparam add_3641_7.INIT0 = 16'h6969;
    defparam add_3641_7.INIT1 = 16'h6969;
    defparam add_3641_7.INJECT1_0 = "NO";
    defparam add_3641_7.INJECT1_1 = "NO";
    CCU2D add_3641_5 (.A0(\B_int[3] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][4] ), 
          .D1(GND_net), .CIN(n62246), .COUT(n62247), .S0(\m_cablesIn[22][4] ), 
          .S1(\m_cablesIn[22][5] ));
    defparam add_3641_5.INIT0 = 16'h6969;
    defparam add_3641_5.INIT1 = 16'h6969;
    defparam add_3641_5.INJECT1_0 = "NO";
    defparam add_3641_5.INJECT1_1 = "NO";
    CCU2D add_3641_3 (.A0(\B_int[1] ), .B0(\QQ_in[21][20] ), .C0(\m_cablesIn[21][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[21][20] ), .C1(\m_cablesIn[21][2] ), 
          .D1(GND_net), .CIN(n62245), .COUT(n62246), .S0(\m_cablesIn[22][2] ), 
          .S1(\m_cablesIn[22][3] ));
    defparam add_3641_3.INIT0 = 16'h6969;
    defparam add_3641_3.INIT1 = 16'h6969;
    defparam add_3641_3.INJECT1_0 = "NO";
    defparam add_3641_3.INJECT1_1 = "NO";
    CCU2D add_3641_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[21][20] ), .C1(\frac_div[6] ), .D1(GND_net), 
          .COUT(n62245), .S1(\m_cablesIn[22][1] ));
    defparam add_3641_1.INIT0 = 16'hF000;
    defparam add_3641_1.INIT1 = 16'h6969;
    defparam add_3641_1.INJECT1_0 = "NO";
    defparam add_3641_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U12 
//

module \a_s(24)_U12  (\m_cablesIn[20][23] , \QQ_in[20][19] , GND_net, 
            \m_cablesIn[20][24] , \m_cablesIn[21][24] , \QQ_in[21][20] , 
            \B_int[21] , \m_cablesIn[20][21] , \B_int[22] , \m_cablesIn[20][22] , 
            \m_cablesIn[21][22] , \m_cablesIn[21][23] , \B_int[19] , \m_cablesIn[20][19] , 
            \B_int[20] , \m_cablesIn[20][20] , \m_cablesIn[21][20] , \m_cablesIn[21][21] , 
            \B_int[17] , \m_cablesIn[20][17] , \B_int[18] , \m_cablesIn[20][18] , 
            \m_cablesIn[21][18] , \m_cablesIn[21][19] , \B_int[15] , \m_cablesIn[20][15] , 
            \B_int[16] , \m_cablesIn[20][16] , \m_cablesIn[21][16] , \m_cablesIn[21][17] , 
            \B_int[13] , \m_cablesIn[20][13] , \B_int[14] , \m_cablesIn[20][14] , 
            \m_cablesIn[21][14] , \m_cablesIn[21][15] , \B_int[11] , \m_cablesIn[20][11] , 
            \B_int[12] , \m_cablesIn[20][12] , \m_cablesIn[21][12] , \m_cablesIn[21][13] , 
            \B_int[9] , \m_cablesIn[20][9] , \B_int[10] , \m_cablesIn[20][10] , 
            \m_cablesIn[21][10] , \m_cablesIn[21][11] , \B_int[7] , \m_cablesIn[20][7] , 
            \B_int[8] , \m_cablesIn[20][8] , \m_cablesIn[21][8] , \m_cablesIn[21][9] , 
            \B_int[5] , \m_cablesIn[20][5] , \B_int[6] , \m_cablesIn[20][6] , 
            \m_cablesIn[21][6] , \m_cablesIn[21][7] , \B_int[3] , \m_cablesIn[20][3] , 
            \B_int[4] , \m_cablesIn[20][4] , \m_cablesIn[21][4] , \m_cablesIn[21][5] , 
            \B_int[1] , \m_cablesIn[20][1] , \B_int[2] , \m_cablesIn[20][2] , 
            \m_cablesIn[21][2] , \m_cablesIn[21][3] , \B_int[0] , \frac_div[7] , 
            \m_cablesIn[21][1] );
    input \m_cablesIn[20][23] ;
    input \QQ_in[20][19] ;
    input GND_net;
    input \m_cablesIn[20][24] ;
    output \m_cablesIn[21][24] ;
    output \QQ_in[21][20] ;
    input \B_int[21] ;
    input \m_cablesIn[20][21] ;
    input \B_int[22] ;
    input \m_cablesIn[20][22] ;
    output \m_cablesIn[21][22] ;
    output \m_cablesIn[21][23] ;
    input \B_int[19] ;
    input \m_cablesIn[20][19] ;
    input \B_int[20] ;
    input \m_cablesIn[20][20] ;
    output \m_cablesIn[21][20] ;
    output \m_cablesIn[21][21] ;
    input \B_int[17] ;
    input \m_cablesIn[20][17] ;
    input \B_int[18] ;
    input \m_cablesIn[20][18] ;
    output \m_cablesIn[21][18] ;
    output \m_cablesIn[21][19] ;
    input \B_int[15] ;
    input \m_cablesIn[20][15] ;
    input \B_int[16] ;
    input \m_cablesIn[20][16] ;
    output \m_cablesIn[21][16] ;
    output \m_cablesIn[21][17] ;
    input \B_int[13] ;
    input \m_cablesIn[20][13] ;
    input \B_int[14] ;
    input \m_cablesIn[20][14] ;
    output \m_cablesIn[21][14] ;
    output \m_cablesIn[21][15] ;
    input \B_int[11] ;
    input \m_cablesIn[20][11] ;
    input \B_int[12] ;
    input \m_cablesIn[20][12] ;
    output \m_cablesIn[21][12] ;
    output \m_cablesIn[21][13] ;
    input \B_int[9] ;
    input \m_cablesIn[20][9] ;
    input \B_int[10] ;
    input \m_cablesIn[20][10] ;
    output \m_cablesIn[21][10] ;
    output \m_cablesIn[21][11] ;
    input \B_int[7] ;
    input \m_cablesIn[20][7] ;
    input \B_int[8] ;
    input \m_cablesIn[20][8] ;
    output \m_cablesIn[21][8] ;
    output \m_cablesIn[21][9] ;
    input \B_int[5] ;
    input \m_cablesIn[20][5] ;
    input \B_int[6] ;
    input \m_cablesIn[20][6] ;
    output \m_cablesIn[21][6] ;
    output \m_cablesIn[21][7] ;
    input \B_int[3] ;
    input \m_cablesIn[20][3] ;
    input \B_int[4] ;
    input \m_cablesIn[20][4] ;
    output \m_cablesIn[21][4] ;
    output \m_cablesIn[21][5] ;
    input \B_int[1] ;
    input \m_cablesIn[20][1] ;
    input \B_int[2] ;
    input \m_cablesIn[20][2] ;
    output \m_cablesIn[21][2] ;
    output \m_cablesIn[21][3] ;
    input \B_int[0] ;
    input \frac_div[7] ;
    output \m_cablesIn[21][1] ;
    
    
    wire n62269, n62268, n62267, n62266, n62265, n62264, n62263, 
        n62262, n62261, n62260, n62259, n62258;
    
    CCU2D add_3615_25 (.A0(\m_cablesIn[20][23] ), .B0(\QQ_in[20][19] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[20][24] ), .B1(\QQ_in[20][19] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62269), .S0(\m_cablesIn[21][24] ), 
          .S1(\QQ_in[21][20] ));
    defparam add_3615_25.INIT0 = 16'h5666;
    defparam add_3615_25.INIT1 = 16'h5999;
    defparam add_3615_25.INJECT1_0 = "NO";
    defparam add_3615_25.INJECT1_1 = "NO";
    CCU2D add_3615_23 (.A0(\B_int[21] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][22] ), 
          .D1(GND_net), .CIN(n62268), .COUT(n62269), .S0(\m_cablesIn[21][22] ), 
          .S1(\m_cablesIn[21][23] ));
    defparam add_3615_23.INIT0 = 16'h6969;
    defparam add_3615_23.INIT1 = 16'h6969;
    defparam add_3615_23.INJECT1_0 = "NO";
    defparam add_3615_23.INJECT1_1 = "NO";
    CCU2D add_3615_21 (.A0(\B_int[19] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][20] ), 
          .D1(GND_net), .CIN(n62267), .COUT(n62268), .S0(\m_cablesIn[21][20] ), 
          .S1(\m_cablesIn[21][21] ));
    defparam add_3615_21.INIT0 = 16'h6969;
    defparam add_3615_21.INIT1 = 16'h6969;
    defparam add_3615_21.INJECT1_0 = "NO";
    defparam add_3615_21.INJECT1_1 = "NO";
    CCU2D add_3615_19 (.A0(\B_int[17] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][18] ), 
          .D1(GND_net), .CIN(n62266), .COUT(n62267), .S0(\m_cablesIn[21][18] ), 
          .S1(\m_cablesIn[21][19] ));
    defparam add_3615_19.INIT0 = 16'h6969;
    defparam add_3615_19.INIT1 = 16'h6969;
    defparam add_3615_19.INJECT1_0 = "NO";
    defparam add_3615_19.INJECT1_1 = "NO";
    CCU2D add_3615_17 (.A0(\B_int[15] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][16] ), 
          .D1(GND_net), .CIN(n62265), .COUT(n62266), .S0(\m_cablesIn[21][16] ), 
          .S1(\m_cablesIn[21][17] ));
    defparam add_3615_17.INIT0 = 16'h6969;
    defparam add_3615_17.INIT1 = 16'h6969;
    defparam add_3615_17.INJECT1_0 = "NO";
    defparam add_3615_17.INJECT1_1 = "NO";
    CCU2D add_3615_15 (.A0(\B_int[13] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][14] ), 
          .D1(GND_net), .CIN(n62264), .COUT(n62265), .S0(\m_cablesIn[21][14] ), 
          .S1(\m_cablesIn[21][15] ));
    defparam add_3615_15.INIT0 = 16'h6969;
    defparam add_3615_15.INIT1 = 16'h6969;
    defparam add_3615_15.INJECT1_0 = "NO";
    defparam add_3615_15.INJECT1_1 = "NO";
    CCU2D add_3615_13 (.A0(\B_int[11] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][12] ), 
          .D1(GND_net), .CIN(n62263), .COUT(n62264), .S0(\m_cablesIn[21][12] ), 
          .S1(\m_cablesIn[21][13] ));
    defparam add_3615_13.INIT0 = 16'h6969;
    defparam add_3615_13.INIT1 = 16'h6969;
    defparam add_3615_13.INJECT1_0 = "NO";
    defparam add_3615_13.INJECT1_1 = "NO";
    CCU2D add_3615_11 (.A0(\B_int[9] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][10] ), 
          .D1(GND_net), .CIN(n62262), .COUT(n62263), .S0(\m_cablesIn[21][10] ), 
          .S1(\m_cablesIn[21][11] ));
    defparam add_3615_11.INIT0 = 16'h6969;
    defparam add_3615_11.INIT1 = 16'h6969;
    defparam add_3615_11.INJECT1_0 = "NO";
    defparam add_3615_11.INJECT1_1 = "NO";
    CCU2D add_3615_9 (.A0(\B_int[7] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][8] ), 
          .D1(GND_net), .CIN(n62261), .COUT(n62262), .S0(\m_cablesIn[21][8] ), 
          .S1(\m_cablesIn[21][9] ));
    defparam add_3615_9.INIT0 = 16'h6969;
    defparam add_3615_9.INIT1 = 16'h6969;
    defparam add_3615_9.INJECT1_0 = "NO";
    defparam add_3615_9.INJECT1_1 = "NO";
    CCU2D add_3615_7 (.A0(\B_int[5] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][6] ), 
          .D1(GND_net), .CIN(n62260), .COUT(n62261), .S0(\m_cablesIn[21][6] ), 
          .S1(\m_cablesIn[21][7] ));
    defparam add_3615_7.INIT0 = 16'h6969;
    defparam add_3615_7.INIT1 = 16'h6969;
    defparam add_3615_7.INJECT1_0 = "NO";
    defparam add_3615_7.INJECT1_1 = "NO";
    CCU2D add_3615_5 (.A0(\B_int[3] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][4] ), 
          .D1(GND_net), .CIN(n62259), .COUT(n62260), .S0(\m_cablesIn[21][4] ), 
          .S1(\m_cablesIn[21][5] ));
    defparam add_3615_5.INIT0 = 16'h6969;
    defparam add_3615_5.INIT1 = 16'h6969;
    defparam add_3615_5.INJECT1_0 = "NO";
    defparam add_3615_5.INJECT1_1 = "NO";
    CCU2D add_3615_3 (.A0(\B_int[1] ), .B0(\QQ_in[20][19] ), .C0(\m_cablesIn[20][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[20][19] ), .C1(\m_cablesIn[20][2] ), 
          .D1(GND_net), .CIN(n62258), .COUT(n62259), .S0(\m_cablesIn[21][2] ), 
          .S1(\m_cablesIn[21][3] ));
    defparam add_3615_3.INIT0 = 16'h6969;
    defparam add_3615_3.INIT1 = 16'h6969;
    defparam add_3615_3.INJECT1_0 = "NO";
    defparam add_3615_3.INJECT1_1 = "NO";
    CCU2D add_3615_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[20][19] ), .C1(\frac_div[7] ), .D1(GND_net), 
          .COUT(n62258), .S1(\m_cablesIn[21][1] ));
    defparam add_3615_1.INIT0 = 16'hF000;
    defparam add_3615_1.INIT1 = 16'h6969;
    defparam add_3615_1.INJECT1_0 = "NO";
    defparam add_3615_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U13 
//

module \a_s(24)_U13  (\m_cablesIn[19][23] , \QQ_in[19][18] , GND_net, 
            \m_cablesIn[19][24] , \m_cablesIn[20][24] , \QQ_in[20][19] , 
            \B_int[21] , \m_cablesIn[19][21] , \B_int[22] , \m_cablesIn[19][22] , 
            \m_cablesIn[20][22] , \m_cablesIn[20][23] , \B_int[19] , \m_cablesIn[19][19] , 
            \B_int[20] , \m_cablesIn[19][20] , \m_cablesIn[20][20] , \m_cablesIn[20][21] , 
            \B_int[17] , \m_cablesIn[19][17] , \B_int[18] , \m_cablesIn[19][18] , 
            \m_cablesIn[20][18] , \m_cablesIn[20][19] , \B_int[15] , \m_cablesIn[19][15] , 
            \B_int[16] , \m_cablesIn[19][16] , \m_cablesIn[20][16] , \m_cablesIn[20][17] , 
            \B_int[13] , \m_cablesIn[19][13] , \B_int[14] , \m_cablesIn[19][14] , 
            \m_cablesIn[20][14] , \m_cablesIn[20][15] , \B_int[11] , \m_cablesIn[19][11] , 
            \B_int[12] , \m_cablesIn[19][12] , \m_cablesIn[20][12] , \m_cablesIn[20][13] , 
            \B_int[9] , \m_cablesIn[19][9] , \B_int[10] , \m_cablesIn[19][10] , 
            \m_cablesIn[20][10] , \m_cablesIn[20][11] , \B_int[7] , \m_cablesIn[19][7] , 
            \B_int[8] , \m_cablesIn[19][8] , \m_cablesIn[20][8] , \m_cablesIn[20][9] , 
            \B_int[5] , \m_cablesIn[19][5] , \B_int[6] , \m_cablesIn[19][6] , 
            \m_cablesIn[20][6] , \m_cablesIn[20][7] , \B_int[3] , \m_cablesIn[19][3] , 
            \B_int[4] , \m_cablesIn[19][4] , \m_cablesIn[20][4] , \m_cablesIn[20][5] , 
            \B_int[1] , \m_cablesIn[19][1] , \B_int[2] , \m_cablesIn[19][2] , 
            \m_cablesIn[20][2] , \m_cablesIn[20][3] , \B_int[0] , \frac_div[8] , 
            \m_cablesIn[20][1] );
    input \m_cablesIn[19][23] ;
    input \QQ_in[19][18] ;
    input GND_net;
    input \m_cablesIn[19][24] ;
    output \m_cablesIn[20][24] ;
    output \QQ_in[20][19] ;
    input \B_int[21] ;
    input \m_cablesIn[19][21] ;
    input \B_int[22] ;
    input \m_cablesIn[19][22] ;
    output \m_cablesIn[20][22] ;
    output \m_cablesIn[20][23] ;
    input \B_int[19] ;
    input \m_cablesIn[19][19] ;
    input \B_int[20] ;
    input \m_cablesIn[19][20] ;
    output \m_cablesIn[20][20] ;
    output \m_cablesIn[20][21] ;
    input \B_int[17] ;
    input \m_cablesIn[19][17] ;
    input \B_int[18] ;
    input \m_cablesIn[19][18] ;
    output \m_cablesIn[20][18] ;
    output \m_cablesIn[20][19] ;
    input \B_int[15] ;
    input \m_cablesIn[19][15] ;
    input \B_int[16] ;
    input \m_cablesIn[19][16] ;
    output \m_cablesIn[20][16] ;
    output \m_cablesIn[20][17] ;
    input \B_int[13] ;
    input \m_cablesIn[19][13] ;
    input \B_int[14] ;
    input \m_cablesIn[19][14] ;
    output \m_cablesIn[20][14] ;
    output \m_cablesIn[20][15] ;
    input \B_int[11] ;
    input \m_cablesIn[19][11] ;
    input \B_int[12] ;
    input \m_cablesIn[19][12] ;
    output \m_cablesIn[20][12] ;
    output \m_cablesIn[20][13] ;
    input \B_int[9] ;
    input \m_cablesIn[19][9] ;
    input \B_int[10] ;
    input \m_cablesIn[19][10] ;
    output \m_cablesIn[20][10] ;
    output \m_cablesIn[20][11] ;
    input \B_int[7] ;
    input \m_cablesIn[19][7] ;
    input \B_int[8] ;
    input \m_cablesIn[19][8] ;
    output \m_cablesIn[20][8] ;
    output \m_cablesIn[20][9] ;
    input \B_int[5] ;
    input \m_cablesIn[19][5] ;
    input \B_int[6] ;
    input \m_cablesIn[19][6] ;
    output \m_cablesIn[20][6] ;
    output \m_cablesIn[20][7] ;
    input \B_int[3] ;
    input \m_cablesIn[19][3] ;
    input \B_int[4] ;
    input \m_cablesIn[19][4] ;
    output \m_cablesIn[20][4] ;
    output \m_cablesIn[20][5] ;
    input \B_int[1] ;
    input \m_cablesIn[19][1] ;
    input \B_int[2] ;
    input \m_cablesIn[19][2] ;
    output \m_cablesIn[20][2] ;
    output \m_cablesIn[20][3] ;
    input \B_int[0] ;
    input \frac_div[8] ;
    output \m_cablesIn[20][1] ;
    
    
    wire n62282, n62281, n62280, n62279, n62278, n62277, n62276, 
        n62275, n62274, n62273, n62272, n62271;
    
    CCU2D add_3589_25 (.A0(\m_cablesIn[19][23] ), .B0(\QQ_in[19][18] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[19][24] ), .B1(\QQ_in[19][18] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62282), .S0(\m_cablesIn[20][24] ), 
          .S1(\QQ_in[20][19] ));
    defparam add_3589_25.INIT0 = 16'h5666;
    defparam add_3589_25.INIT1 = 16'h5999;
    defparam add_3589_25.INJECT1_0 = "NO";
    defparam add_3589_25.INJECT1_1 = "NO";
    CCU2D add_3589_23 (.A0(\B_int[21] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][22] ), 
          .D1(GND_net), .CIN(n62281), .COUT(n62282), .S0(\m_cablesIn[20][22] ), 
          .S1(\m_cablesIn[20][23] ));
    defparam add_3589_23.INIT0 = 16'h6969;
    defparam add_3589_23.INIT1 = 16'h6969;
    defparam add_3589_23.INJECT1_0 = "NO";
    defparam add_3589_23.INJECT1_1 = "NO";
    CCU2D add_3589_21 (.A0(\B_int[19] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][20] ), 
          .D1(GND_net), .CIN(n62280), .COUT(n62281), .S0(\m_cablesIn[20][20] ), 
          .S1(\m_cablesIn[20][21] ));
    defparam add_3589_21.INIT0 = 16'h6969;
    defparam add_3589_21.INIT1 = 16'h6969;
    defparam add_3589_21.INJECT1_0 = "NO";
    defparam add_3589_21.INJECT1_1 = "NO";
    CCU2D add_3589_19 (.A0(\B_int[17] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][18] ), 
          .D1(GND_net), .CIN(n62279), .COUT(n62280), .S0(\m_cablesIn[20][18] ), 
          .S1(\m_cablesIn[20][19] ));
    defparam add_3589_19.INIT0 = 16'h6969;
    defparam add_3589_19.INIT1 = 16'h6969;
    defparam add_3589_19.INJECT1_0 = "NO";
    defparam add_3589_19.INJECT1_1 = "NO";
    CCU2D add_3589_17 (.A0(\B_int[15] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][16] ), 
          .D1(GND_net), .CIN(n62278), .COUT(n62279), .S0(\m_cablesIn[20][16] ), 
          .S1(\m_cablesIn[20][17] ));
    defparam add_3589_17.INIT0 = 16'h6969;
    defparam add_3589_17.INIT1 = 16'h6969;
    defparam add_3589_17.INJECT1_0 = "NO";
    defparam add_3589_17.INJECT1_1 = "NO";
    CCU2D add_3589_15 (.A0(\B_int[13] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][14] ), 
          .D1(GND_net), .CIN(n62277), .COUT(n62278), .S0(\m_cablesIn[20][14] ), 
          .S1(\m_cablesIn[20][15] ));
    defparam add_3589_15.INIT0 = 16'h6969;
    defparam add_3589_15.INIT1 = 16'h6969;
    defparam add_3589_15.INJECT1_0 = "NO";
    defparam add_3589_15.INJECT1_1 = "NO";
    CCU2D add_3589_13 (.A0(\B_int[11] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][12] ), 
          .D1(GND_net), .CIN(n62276), .COUT(n62277), .S0(\m_cablesIn[20][12] ), 
          .S1(\m_cablesIn[20][13] ));
    defparam add_3589_13.INIT0 = 16'h6969;
    defparam add_3589_13.INIT1 = 16'h6969;
    defparam add_3589_13.INJECT1_0 = "NO";
    defparam add_3589_13.INJECT1_1 = "NO";
    CCU2D add_3589_11 (.A0(\B_int[9] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][10] ), 
          .D1(GND_net), .CIN(n62275), .COUT(n62276), .S0(\m_cablesIn[20][10] ), 
          .S1(\m_cablesIn[20][11] ));
    defparam add_3589_11.INIT0 = 16'h6969;
    defparam add_3589_11.INIT1 = 16'h6969;
    defparam add_3589_11.INJECT1_0 = "NO";
    defparam add_3589_11.INJECT1_1 = "NO";
    CCU2D add_3589_9 (.A0(\B_int[7] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][8] ), 
          .D1(GND_net), .CIN(n62274), .COUT(n62275), .S0(\m_cablesIn[20][8] ), 
          .S1(\m_cablesIn[20][9] ));
    defparam add_3589_9.INIT0 = 16'h6969;
    defparam add_3589_9.INIT1 = 16'h6969;
    defparam add_3589_9.INJECT1_0 = "NO";
    defparam add_3589_9.INJECT1_1 = "NO";
    CCU2D add_3589_7 (.A0(\B_int[5] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][6] ), 
          .D1(GND_net), .CIN(n62273), .COUT(n62274), .S0(\m_cablesIn[20][6] ), 
          .S1(\m_cablesIn[20][7] ));
    defparam add_3589_7.INIT0 = 16'h6969;
    defparam add_3589_7.INIT1 = 16'h6969;
    defparam add_3589_7.INJECT1_0 = "NO";
    defparam add_3589_7.INJECT1_1 = "NO";
    CCU2D add_3589_5 (.A0(\B_int[3] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][4] ), 
          .D1(GND_net), .CIN(n62272), .COUT(n62273), .S0(\m_cablesIn[20][4] ), 
          .S1(\m_cablesIn[20][5] ));
    defparam add_3589_5.INIT0 = 16'h6969;
    defparam add_3589_5.INIT1 = 16'h6969;
    defparam add_3589_5.INJECT1_0 = "NO";
    defparam add_3589_5.INJECT1_1 = "NO";
    CCU2D add_3589_3 (.A0(\B_int[1] ), .B0(\QQ_in[19][18] ), .C0(\m_cablesIn[19][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[19][18] ), .C1(\m_cablesIn[19][2] ), 
          .D1(GND_net), .CIN(n62271), .COUT(n62272), .S0(\m_cablesIn[20][2] ), 
          .S1(\m_cablesIn[20][3] ));
    defparam add_3589_3.INIT0 = 16'h6969;
    defparam add_3589_3.INIT1 = 16'h6969;
    defparam add_3589_3.INJECT1_0 = "NO";
    defparam add_3589_3.INJECT1_1 = "NO";
    CCU2D add_3589_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[19][18] ), .C1(\frac_div[8] ), .D1(GND_net), 
          .COUT(n62271), .S1(\m_cablesIn[20][1] ));
    defparam add_3589_1.INIT0 = 16'hF000;
    defparam add_3589_1.INIT1 = 16'h6969;
    defparam add_3589_1.INJECT1_0 = "NO";
    defparam add_3589_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U14 
//

module \a_s(24)_U14  (GND_net, \m_cablesIn[1][24] , \QQ_in[1][0] , \A_int[21] , 
            \B_int[21] , \A_int[22] , \B_int[22] , \m_cablesIn[1][22] , 
            \m_cablesIn[1][23] , \A_int[19] , \B_int[19] , \A_int[20] , 
            \B_int[20] , \m_cablesIn[1][20] , \m_cablesIn[1][21] , \A_int[17] , 
            \B_int[17] , \A_int[18] , \B_int[18] , \m_cablesIn[1][18] , 
            \m_cablesIn[1][19] , \A_int[15] , \B_int[15] , \A_int[16] , 
            \B_int[16] , \m_cablesIn[1][16] , \m_cablesIn[1][17] , \A_int[13] , 
            \B_int[13] , \A_int[14] , \B_int[14] , \m_cablesIn[1][14] , 
            \m_cablesIn[1][15] , \A_int[11] , \B_int[11] , \A_int[12] , 
            \B_int[12] , \m_cablesIn[1][12] , \m_cablesIn[1][13] , \A_int[9] , 
            \B_int[9] , \A_int[10] , \B_int[10] , \m_cablesIn[1][10] , 
            \m_cablesIn[1][11] , \A_int[7] , \B_int[7] , \A_int[8] , 
            \B_int[8] , \m_cablesIn[1][8] , \m_cablesIn[1][9] , \A_int[5] , 
            \B_int[5] , \A_int[6] , \B_int[6] , \m_cablesIn[1][6] , 
            \m_cablesIn[1][7] , \A_int[3] , \B_int[3] , \A_int[4] , 
            \B_int[4] , \m_cablesIn[1][4] , \m_cablesIn[1][5] , \A_int[1] , 
            \B_int[1] , \A_int[2] , \B_int[2] , \m_cablesIn[1][2] , 
            \m_cablesIn[1][3] , \A_int[0] , \B_int[0] , \m_cablesIn[1][1] );
    input GND_net;
    output \m_cablesIn[1][24] ;
    output \QQ_in[1][0] ;
    input \A_int[21] ;
    input \B_int[21] ;
    input \A_int[22] ;
    input \B_int[22] ;
    output \m_cablesIn[1][22] ;
    output \m_cablesIn[1][23] ;
    input \A_int[19] ;
    input \B_int[19] ;
    input \A_int[20] ;
    input \B_int[20] ;
    output \m_cablesIn[1][20] ;
    output \m_cablesIn[1][21] ;
    input \A_int[17] ;
    input \B_int[17] ;
    input \A_int[18] ;
    input \B_int[18] ;
    output \m_cablesIn[1][18] ;
    output \m_cablesIn[1][19] ;
    input \A_int[15] ;
    input \B_int[15] ;
    input \A_int[16] ;
    input \B_int[16] ;
    output \m_cablesIn[1][16] ;
    output \m_cablesIn[1][17] ;
    input \A_int[13] ;
    input \B_int[13] ;
    input \A_int[14] ;
    input \B_int[14] ;
    output \m_cablesIn[1][14] ;
    output \m_cablesIn[1][15] ;
    input \A_int[11] ;
    input \B_int[11] ;
    input \A_int[12] ;
    input \B_int[12] ;
    output \m_cablesIn[1][12] ;
    output \m_cablesIn[1][13] ;
    input \A_int[9] ;
    input \B_int[9] ;
    input \A_int[10] ;
    input \B_int[10] ;
    output \m_cablesIn[1][10] ;
    output \m_cablesIn[1][11] ;
    input \A_int[7] ;
    input \B_int[7] ;
    input \A_int[8] ;
    input \B_int[8] ;
    output \m_cablesIn[1][8] ;
    output \m_cablesIn[1][9] ;
    input \A_int[5] ;
    input \B_int[5] ;
    input \A_int[6] ;
    input \B_int[6] ;
    output \m_cablesIn[1][6] ;
    output \m_cablesIn[1][7] ;
    input \A_int[3] ;
    input \B_int[3] ;
    input \A_int[4] ;
    input \B_int[4] ;
    output \m_cablesIn[1][4] ;
    output \m_cablesIn[1][5] ;
    input \A_int[1] ;
    input \B_int[1] ;
    input \A_int[2] ;
    input \B_int[2] ;
    output \m_cablesIn[1][2] ;
    output \m_cablesIn[1][3] ;
    input \A_int[0] ;
    input \B_int[0] ;
    output \m_cablesIn[1][1] ;
    
    
    wire n62167, n62166, n62165, n62164, n62163, n62162, n62161, 
        n62160, n62159, n62158, n62157, n62156;
    
    CCU2D sub_8_add_2_25 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62167), 
          .S0(\m_cablesIn[1][24] ), .S1(\QQ_in[1][0] ));
    defparam sub_8_add_2_25.INIT0 = 16'h0fff;
    defparam sub_8_add_2_25.INIT1 = 16'hffff;
    defparam sub_8_add_2_25.INJECT1_0 = "NO";
    defparam sub_8_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_23 (.A0(\A_int[21] ), .B0(\B_int[21] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[22] ), .B1(\B_int[22] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62166), .COUT(n62167), .S0(\m_cablesIn[1][22] ), 
          .S1(\m_cablesIn[1][23] ));
    defparam sub_8_add_2_23.INIT0 = 16'h5999;
    defparam sub_8_add_2_23.INIT1 = 16'h5999;
    defparam sub_8_add_2_23.INJECT1_0 = "NO";
    defparam sub_8_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_21 (.A0(\A_int[19] ), .B0(\B_int[19] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[20] ), .B1(\B_int[20] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62165), .COUT(n62166), .S0(\m_cablesIn[1][20] ), 
          .S1(\m_cablesIn[1][21] ));
    defparam sub_8_add_2_21.INIT0 = 16'h5999;
    defparam sub_8_add_2_21.INIT1 = 16'h5999;
    defparam sub_8_add_2_21.INJECT1_0 = "NO";
    defparam sub_8_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_19 (.A0(\A_int[17] ), .B0(\B_int[17] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[18] ), .B1(\B_int[18] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62164), .COUT(n62165), .S0(\m_cablesIn[1][18] ), 
          .S1(\m_cablesIn[1][19] ));
    defparam sub_8_add_2_19.INIT0 = 16'h5999;
    defparam sub_8_add_2_19.INIT1 = 16'h5999;
    defparam sub_8_add_2_19.INJECT1_0 = "NO";
    defparam sub_8_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_17 (.A0(\A_int[15] ), .B0(\B_int[15] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[16] ), .B1(\B_int[16] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62163), .COUT(n62164), .S0(\m_cablesIn[1][16] ), 
          .S1(\m_cablesIn[1][17] ));
    defparam sub_8_add_2_17.INIT0 = 16'h5999;
    defparam sub_8_add_2_17.INIT1 = 16'h5999;
    defparam sub_8_add_2_17.INJECT1_0 = "NO";
    defparam sub_8_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_15 (.A0(\A_int[13] ), .B0(\B_int[13] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[14] ), .B1(\B_int[14] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62162), .COUT(n62163), .S0(\m_cablesIn[1][14] ), 
          .S1(\m_cablesIn[1][15] ));
    defparam sub_8_add_2_15.INIT0 = 16'h5999;
    defparam sub_8_add_2_15.INIT1 = 16'h5999;
    defparam sub_8_add_2_15.INJECT1_0 = "NO";
    defparam sub_8_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_13 (.A0(\A_int[11] ), .B0(\B_int[11] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[12] ), .B1(\B_int[12] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62161), .COUT(n62162), .S0(\m_cablesIn[1][12] ), 
          .S1(\m_cablesIn[1][13] ));
    defparam sub_8_add_2_13.INIT0 = 16'h5999;
    defparam sub_8_add_2_13.INIT1 = 16'h5999;
    defparam sub_8_add_2_13.INJECT1_0 = "NO";
    defparam sub_8_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_11 (.A0(\A_int[9] ), .B0(\B_int[9] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[10] ), .B1(\B_int[10] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62160), .COUT(n62161), .S0(\m_cablesIn[1][10] ), 
          .S1(\m_cablesIn[1][11] ));
    defparam sub_8_add_2_11.INIT0 = 16'h5999;
    defparam sub_8_add_2_11.INIT1 = 16'h5999;
    defparam sub_8_add_2_11.INJECT1_0 = "NO";
    defparam sub_8_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_9 (.A0(\A_int[7] ), .B0(\B_int[7] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[8] ), .B1(\B_int[8] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62159), .COUT(n62160), .S0(\m_cablesIn[1][8] ), 
          .S1(\m_cablesIn[1][9] ));
    defparam sub_8_add_2_9.INIT0 = 16'h5999;
    defparam sub_8_add_2_9.INIT1 = 16'h5999;
    defparam sub_8_add_2_9.INJECT1_0 = "NO";
    defparam sub_8_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_7 (.A0(\A_int[5] ), .B0(\B_int[5] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[6] ), .B1(\B_int[6] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62158), .COUT(n62159), .S0(\m_cablesIn[1][6] ), 
          .S1(\m_cablesIn[1][7] ));
    defparam sub_8_add_2_7.INIT0 = 16'h5999;
    defparam sub_8_add_2_7.INIT1 = 16'h5999;
    defparam sub_8_add_2_7.INJECT1_0 = "NO";
    defparam sub_8_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_5 (.A0(\A_int[3] ), .B0(\B_int[3] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[4] ), .B1(\B_int[4] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62157), .COUT(n62158), .S0(\m_cablesIn[1][4] ), 
          .S1(\m_cablesIn[1][5] ));
    defparam sub_8_add_2_5.INIT0 = 16'h5999;
    defparam sub_8_add_2_5.INIT1 = 16'h5999;
    defparam sub_8_add_2_5.INJECT1_0 = "NO";
    defparam sub_8_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_3 (.A0(\A_int[1] ), .B0(\B_int[1] ), .C0(GND_net), 
          .D0(GND_net), .A1(\A_int[2] ), .B1(\B_int[2] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n62156), .COUT(n62157), .S0(\m_cablesIn[1][2] ), 
          .S1(\m_cablesIn[1][3] ));
    defparam sub_8_add_2_3.INIT0 = 16'h5999;
    defparam sub_8_add_2_3.INIT1 = 16'h5999;
    defparam sub_8_add_2_3.INJECT1_0 = "NO";
    defparam sub_8_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\A_int[0] ), .B1(\B_int[0] ), .C1(GND_net), .D1(GND_net), 
          .COUT(n62156), .S1(\m_cablesIn[1][1] ));
    defparam sub_8_add_2_1.INIT0 = 16'h0000;
    defparam sub_8_add_2_1.INIT1 = 16'h5999;
    defparam sub_8_add_2_1.INJECT1_0 = "NO";
    defparam sub_8_add_2_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U15 
//

module \a_s(24)_U15  (\m_cablesIn[18][23] , \QQ_in[18][17] , GND_net, 
            \m_cablesIn[18][24] , \m_cablesIn[19][24] , \QQ_in[19][18] , 
            \B_int[21] , \m_cablesIn[18][21] , \B_int[22] , \m_cablesIn[18][22] , 
            \m_cablesIn[19][22] , \m_cablesIn[19][23] , \B_int[19] , \m_cablesIn[18][19] , 
            \B_int[20] , \m_cablesIn[18][20] , \m_cablesIn[19][20] , \m_cablesIn[19][21] , 
            \B_int[17] , \m_cablesIn[18][17] , \B_int[18] , \m_cablesIn[18][18] , 
            \m_cablesIn[19][18] , \m_cablesIn[19][19] , \B_int[15] , \m_cablesIn[18][15] , 
            \B_int[16] , \m_cablesIn[18][16] , \m_cablesIn[19][16] , \m_cablesIn[19][17] , 
            \B_int[13] , \m_cablesIn[18][13] , \B_int[14] , \m_cablesIn[18][14] , 
            \m_cablesIn[19][14] , \m_cablesIn[19][15] , \B_int[11] , \m_cablesIn[18][11] , 
            \B_int[12] , \m_cablesIn[18][12] , \m_cablesIn[19][12] , \m_cablesIn[19][13] , 
            \B_int[9] , \m_cablesIn[18][9] , \B_int[10] , \m_cablesIn[18][10] , 
            \m_cablesIn[19][10] , \m_cablesIn[19][11] , \B_int[7] , \m_cablesIn[18][7] , 
            \B_int[8] , \m_cablesIn[18][8] , \m_cablesIn[19][8] , \m_cablesIn[19][9] , 
            \B_int[5] , \m_cablesIn[18][5] , \B_int[6] , \m_cablesIn[18][6] , 
            \m_cablesIn[19][6] , \m_cablesIn[19][7] , \B_int[3] , \m_cablesIn[18][3] , 
            \B_int[4] , \m_cablesIn[18][4] , \m_cablesIn[19][4] , \m_cablesIn[19][5] , 
            \B_int[1] , \m_cablesIn[18][1] , \B_int[2] , \m_cablesIn[18][2] , 
            \m_cablesIn[19][2] , \m_cablesIn[19][3] , \B_int[0] , \frac_div[9] , 
            \m_cablesIn[19][1] );
    input \m_cablesIn[18][23] ;
    input \QQ_in[18][17] ;
    input GND_net;
    input \m_cablesIn[18][24] ;
    output \m_cablesIn[19][24] ;
    output \QQ_in[19][18] ;
    input \B_int[21] ;
    input \m_cablesIn[18][21] ;
    input \B_int[22] ;
    input \m_cablesIn[18][22] ;
    output \m_cablesIn[19][22] ;
    output \m_cablesIn[19][23] ;
    input \B_int[19] ;
    input \m_cablesIn[18][19] ;
    input \B_int[20] ;
    input \m_cablesIn[18][20] ;
    output \m_cablesIn[19][20] ;
    output \m_cablesIn[19][21] ;
    input \B_int[17] ;
    input \m_cablesIn[18][17] ;
    input \B_int[18] ;
    input \m_cablesIn[18][18] ;
    output \m_cablesIn[19][18] ;
    output \m_cablesIn[19][19] ;
    input \B_int[15] ;
    input \m_cablesIn[18][15] ;
    input \B_int[16] ;
    input \m_cablesIn[18][16] ;
    output \m_cablesIn[19][16] ;
    output \m_cablesIn[19][17] ;
    input \B_int[13] ;
    input \m_cablesIn[18][13] ;
    input \B_int[14] ;
    input \m_cablesIn[18][14] ;
    output \m_cablesIn[19][14] ;
    output \m_cablesIn[19][15] ;
    input \B_int[11] ;
    input \m_cablesIn[18][11] ;
    input \B_int[12] ;
    input \m_cablesIn[18][12] ;
    output \m_cablesIn[19][12] ;
    output \m_cablesIn[19][13] ;
    input \B_int[9] ;
    input \m_cablesIn[18][9] ;
    input \B_int[10] ;
    input \m_cablesIn[18][10] ;
    output \m_cablesIn[19][10] ;
    output \m_cablesIn[19][11] ;
    input \B_int[7] ;
    input \m_cablesIn[18][7] ;
    input \B_int[8] ;
    input \m_cablesIn[18][8] ;
    output \m_cablesIn[19][8] ;
    output \m_cablesIn[19][9] ;
    input \B_int[5] ;
    input \m_cablesIn[18][5] ;
    input \B_int[6] ;
    input \m_cablesIn[18][6] ;
    output \m_cablesIn[19][6] ;
    output \m_cablesIn[19][7] ;
    input \B_int[3] ;
    input \m_cablesIn[18][3] ;
    input \B_int[4] ;
    input \m_cablesIn[18][4] ;
    output \m_cablesIn[19][4] ;
    output \m_cablesIn[19][5] ;
    input \B_int[1] ;
    input \m_cablesIn[18][1] ;
    input \B_int[2] ;
    input \m_cablesIn[18][2] ;
    output \m_cablesIn[19][2] ;
    output \m_cablesIn[19][3] ;
    input \B_int[0] ;
    input \frac_div[9] ;
    output \m_cablesIn[19][1] ;
    
    
    wire n62295, n62294, n62293, n62292, n62291, n62290, n62289, 
        n62288, n62287, n62286, n62285, n62284;
    
    CCU2D add_3563_25 (.A0(\m_cablesIn[18][23] ), .B0(\QQ_in[18][17] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[18][24] ), .B1(\QQ_in[18][17] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62295), .S0(\m_cablesIn[19][24] ), 
          .S1(\QQ_in[19][18] ));
    defparam add_3563_25.INIT0 = 16'h5666;
    defparam add_3563_25.INIT1 = 16'h5999;
    defparam add_3563_25.INJECT1_0 = "NO";
    defparam add_3563_25.INJECT1_1 = "NO";
    CCU2D add_3563_23 (.A0(\B_int[21] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][22] ), 
          .D1(GND_net), .CIN(n62294), .COUT(n62295), .S0(\m_cablesIn[19][22] ), 
          .S1(\m_cablesIn[19][23] ));
    defparam add_3563_23.INIT0 = 16'h6969;
    defparam add_3563_23.INIT1 = 16'h6969;
    defparam add_3563_23.INJECT1_0 = "NO";
    defparam add_3563_23.INJECT1_1 = "NO";
    CCU2D add_3563_21 (.A0(\B_int[19] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][20] ), 
          .D1(GND_net), .CIN(n62293), .COUT(n62294), .S0(\m_cablesIn[19][20] ), 
          .S1(\m_cablesIn[19][21] ));
    defparam add_3563_21.INIT0 = 16'h6969;
    defparam add_3563_21.INIT1 = 16'h6969;
    defparam add_3563_21.INJECT1_0 = "NO";
    defparam add_3563_21.INJECT1_1 = "NO";
    CCU2D add_3563_19 (.A0(\B_int[17] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][18] ), 
          .D1(GND_net), .CIN(n62292), .COUT(n62293), .S0(\m_cablesIn[19][18] ), 
          .S1(\m_cablesIn[19][19] ));
    defparam add_3563_19.INIT0 = 16'h6969;
    defparam add_3563_19.INIT1 = 16'h6969;
    defparam add_3563_19.INJECT1_0 = "NO";
    defparam add_3563_19.INJECT1_1 = "NO";
    CCU2D add_3563_17 (.A0(\B_int[15] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][16] ), 
          .D1(GND_net), .CIN(n62291), .COUT(n62292), .S0(\m_cablesIn[19][16] ), 
          .S1(\m_cablesIn[19][17] ));
    defparam add_3563_17.INIT0 = 16'h6969;
    defparam add_3563_17.INIT1 = 16'h6969;
    defparam add_3563_17.INJECT1_0 = "NO";
    defparam add_3563_17.INJECT1_1 = "NO";
    CCU2D add_3563_15 (.A0(\B_int[13] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][14] ), 
          .D1(GND_net), .CIN(n62290), .COUT(n62291), .S0(\m_cablesIn[19][14] ), 
          .S1(\m_cablesIn[19][15] ));
    defparam add_3563_15.INIT0 = 16'h6969;
    defparam add_3563_15.INIT1 = 16'h6969;
    defparam add_3563_15.INJECT1_0 = "NO";
    defparam add_3563_15.INJECT1_1 = "NO";
    CCU2D add_3563_13 (.A0(\B_int[11] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][12] ), 
          .D1(GND_net), .CIN(n62289), .COUT(n62290), .S0(\m_cablesIn[19][12] ), 
          .S1(\m_cablesIn[19][13] ));
    defparam add_3563_13.INIT0 = 16'h6969;
    defparam add_3563_13.INIT1 = 16'h6969;
    defparam add_3563_13.INJECT1_0 = "NO";
    defparam add_3563_13.INJECT1_1 = "NO";
    CCU2D add_3563_11 (.A0(\B_int[9] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][10] ), 
          .D1(GND_net), .CIN(n62288), .COUT(n62289), .S0(\m_cablesIn[19][10] ), 
          .S1(\m_cablesIn[19][11] ));
    defparam add_3563_11.INIT0 = 16'h6969;
    defparam add_3563_11.INIT1 = 16'h6969;
    defparam add_3563_11.INJECT1_0 = "NO";
    defparam add_3563_11.INJECT1_1 = "NO";
    CCU2D add_3563_9 (.A0(\B_int[7] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][8] ), 
          .D1(GND_net), .CIN(n62287), .COUT(n62288), .S0(\m_cablesIn[19][8] ), 
          .S1(\m_cablesIn[19][9] ));
    defparam add_3563_9.INIT0 = 16'h6969;
    defparam add_3563_9.INIT1 = 16'h6969;
    defparam add_3563_9.INJECT1_0 = "NO";
    defparam add_3563_9.INJECT1_1 = "NO";
    CCU2D add_3563_7 (.A0(\B_int[5] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][6] ), 
          .D1(GND_net), .CIN(n62286), .COUT(n62287), .S0(\m_cablesIn[19][6] ), 
          .S1(\m_cablesIn[19][7] ));
    defparam add_3563_7.INIT0 = 16'h6969;
    defparam add_3563_7.INIT1 = 16'h6969;
    defparam add_3563_7.INJECT1_0 = "NO";
    defparam add_3563_7.INJECT1_1 = "NO";
    CCU2D add_3563_5 (.A0(\B_int[3] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][4] ), 
          .D1(GND_net), .CIN(n62285), .COUT(n62286), .S0(\m_cablesIn[19][4] ), 
          .S1(\m_cablesIn[19][5] ));
    defparam add_3563_5.INIT0 = 16'h6969;
    defparam add_3563_5.INIT1 = 16'h6969;
    defparam add_3563_5.INJECT1_0 = "NO";
    defparam add_3563_5.INJECT1_1 = "NO";
    CCU2D add_3563_3 (.A0(\B_int[1] ), .B0(\QQ_in[18][17] ), .C0(\m_cablesIn[18][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[18][17] ), .C1(\m_cablesIn[18][2] ), 
          .D1(GND_net), .CIN(n62284), .COUT(n62285), .S0(\m_cablesIn[19][2] ), 
          .S1(\m_cablesIn[19][3] ));
    defparam add_3563_3.INIT0 = 16'h6969;
    defparam add_3563_3.INIT1 = 16'h6969;
    defparam add_3563_3.INJECT1_0 = "NO";
    defparam add_3563_3.INJECT1_1 = "NO";
    CCU2D add_3563_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[18][17] ), .C1(\frac_div[9] ), .D1(GND_net), 
          .COUT(n62284), .S1(\m_cablesIn[19][1] ));
    defparam add_3563_1.INIT0 = 16'hF000;
    defparam add_3563_1.INIT1 = 16'h6969;
    defparam add_3563_1.INJECT1_0 = "NO";
    defparam add_3563_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U16 
//

module \a_s(24)_U16  (\m_cablesIn[17][23] , \QQ_in[17][16] , GND_net, 
            \m_cablesIn[17][24] , \m_cablesIn[18][24] , \QQ_in[18][17] , 
            \B_int[21] , \m_cablesIn[17][21] , \B_int[22] , \m_cablesIn[17][22] , 
            \m_cablesIn[18][22] , \m_cablesIn[18][23] , \B_int[19] , \m_cablesIn[17][19] , 
            \B_int[20] , \m_cablesIn[17][20] , \m_cablesIn[18][20] , \m_cablesIn[18][21] , 
            \B_int[17] , \m_cablesIn[17][17] , \B_int[18] , \m_cablesIn[17][18] , 
            \m_cablesIn[18][18] , \m_cablesIn[18][19] , \B_int[15] , \m_cablesIn[17][15] , 
            \B_int[16] , \m_cablesIn[17][16] , \m_cablesIn[18][16] , \m_cablesIn[18][17] , 
            \B_int[13] , \m_cablesIn[17][13] , \B_int[14] , \m_cablesIn[17][14] , 
            \m_cablesIn[18][14] , \m_cablesIn[18][15] , \B_int[11] , \m_cablesIn[17][11] , 
            \B_int[12] , \m_cablesIn[17][12] , \m_cablesIn[18][12] , \m_cablesIn[18][13] , 
            \B_int[9] , \m_cablesIn[17][9] , \B_int[10] , \m_cablesIn[17][10] , 
            \m_cablesIn[18][10] , \m_cablesIn[18][11] , \B_int[7] , \m_cablesIn[17][7] , 
            \B_int[8] , \m_cablesIn[17][8] , \m_cablesIn[18][8] , \m_cablesIn[18][9] , 
            \B_int[5] , \m_cablesIn[17][5] , \B_int[6] , \m_cablesIn[17][6] , 
            \m_cablesIn[18][6] , \m_cablesIn[18][7] , \B_int[3] , \m_cablesIn[17][3] , 
            \B_int[4] , \m_cablesIn[17][4] , \m_cablesIn[18][4] , \m_cablesIn[18][5] , 
            \B_int[1] , \m_cablesIn[17][1] , \B_int[2] , \m_cablesIn[17][2] , 
            \m_cablesIn[18][2] , \m_cablesIn[18][3] , \B_int[0] , \frac_div[10] , 
            \m_cablesIn[18][1] );
    input \m_cablesIn[17][23] ;
    input \QQ_in[17][16] ;
    input GND_net;
    input \m_cablesIn[17][24] ;
    output \m_cablesIn[18][24] ;
    output \QQ_in[18][17] ;
    input \B_int[21] ;
    input \m_cablesIn[17][21] ;
    input \B_int[22] ;
    input \m_cablesIn[17][22] ;
    output \m_cablesIn[18][22] ;
    output \m_cablesIn[18][23] ;
    input \B_int[19] ;
    input \m_cablesIn[17][19] ;
    input \B_int[20] ;
    input \m_cablesIn[17][20] ;
    output \m_cablesIn[18][20] ;
    output \m_cablesIn[18][21] ;
    input \B_int[17] ;
    input \m_cablesIn[17][17] ;
    input \B_int[18] ;
    input \m_cablesIn[17][18] ;
    output \m_cablesIn[18][18] ;
    output \m_cablesIn[18][19] ;
    input \B_int[15] ;
    input \m_cablesIn[17][15] ;
    input \B_int[16] ;
    input \m_cablesIn[17][16] ;
    output \m_cablesIn[18][16] ;
    output \m_cablesIn[18][17] ;
    input \B_int[13] ;
    input \m_cablesIn[17][13] ;
    input \B_int[14] ;
    input \m_cablesIn[17][14] ;
    output \m_cablesIn[18][14] ;
    output \m_cablesIn[18][15] ;
    input \B_int[11] ;
    input \m_cablesIn[17][11] ;
    input \B_int[12] ;
    input \m_cablesIn[17][12] ;
    output \m_cablesIn[18][12] ;
    output \m_cablesIn[18][13] ;
    input \B_int[9] ;
    input \m_cablesIn[17][9] ;
    input \B_int[10] ;
    input \m_cablesIn[17][10] ;
    output \m_cablesIn[18][10] ;
    output \m_cablesIn[18][11] ;
    input \B_int[7] ;
    input \m_cablesIn[17][7] ;
    input \B_int[8] ;
    input \m_cablesIn[17][8] ;
    output \m_cablesIn[18][8] ;
    output \m_cablesIn[18][9] ;
    input \B_int[5] ;
    input \m_cablesIn[17][5] ;
    input \B_int[6] ;
    input \m_cablesIn[17][6] ;
    output \m_cablesIn[18][6] ;
    output \m_cablesIn[18][7] ;
    input \B_int[3] ;
    input \m_cablesIn[17][3] ;
    input \B_int[4] ;
    input \m_cablesIn[17][4] ;
    output \m_cablesIn[18][4] ;
    output \m_cablesIn[18][5] ;
    input \B_int[1] ;
    input \m_cablesIn[17][1] ;
    input \B_int[2] ;
    input \m_cablesIn[17][2] ;
    output \m_cablesIn[18][2] ;
    output \m_cablesIn[18][3] ;
    input \B_int[0] ;
    input \frac_div[10] ;
    output \m_cablesIn[18][1] ;
    
    
    wire n62308, n62307, n62306, n62305, n62304, n62303, n62302, 
        n62301, n62300, n62299, n62298, n62297;
    
    CCU2D add_3537_25 (.A0(\m_cablesIn[17][23] ), .B0(\QQ_in[17][16] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[17][24] ), .B1(\QQ_in[17][16] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62308), .S0(\m_cablesIn[18][24] ), 
          .S1(\QQ_in[18][17] ));
    defparam add_3537_25.INIT0 = 16'h5666;
    defparam add_3537_25.INIT1 = 16'h5999;
    defparam add_3537_25.INJECT1_0 = "NO";
    defparam add_3537_25.INJECT1_1 = "NO";
    CCU2D add_3537_23 (.A0(\B_int[21] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][22] ), 
          .D1(GND_net), .CIN(n62307), .COUT(n62308), .S0(\m_cablesIn[18][22] ), 
          .S1(\m_cablesIn[18][23] ));
    defparam add_3537_23.INIT0 = 16'h6969;
    defparam add_3537_23.INIT1 = 16'h6969;
    defparam add_3537_23.INJECT1_0 = "NO";
    defparam add_3537_23.INJECT1_1 = "NO";
    CCU2D add_3537_21 (.A0(\B_int[19] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][20] ), 
          .D1(GND_net), .CIN(n62306), .COUT(n62307), .S0(\m_cablesIn[18][20] ), 
          .S1(\m_cablesIn[18][21] ));
    defparam add_3537_21.INIT0 = 16'h6969;
    defparam add_3537_21.INIT1 = 16'h6969;
    defparam add_3537_21.INJECT1_0 = "NO";
    defparam add_3537_21.INJECT1_1 = "NO";
    CCU2D add_3537_19 (.A0(\B_int[17] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][18] ), 
          .D1(GND_net), .CIN(n62305), .COUT(n62306), .S0(\m_cablesIn[18][18] ), 
          .S1(\m_cablesIn[18][19] ));
    defparam add_3537_19.INIT0 = 16'h6969;
    defparam add_3537_19.INIT1 = 16'h6969;
    defparam add_3537_19.INJECT1_0 = "NO";
    defparam add_3537_19.INJECT1_1 = "NO";
    CCU2D add_3537_17 (.A0(\B_int[15] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][16] ), 
          .D1(GND_net), .CIN(n62304), .COUT(n62305), .S0(\m_cablesIn[18][16] ), 
          .S1(\m_cablesIn[18][17] ));
    defparam add_3537_17.INIT0 = 16'h6969;
    defparam add_3537_17.INIT1 = 16'h6969;
    defparam add_3537_17.INJECT1_0 = "NO";
    defparam add_3537_17.INJECT1_1 = "NO";
    CCU2D add_3537_15 (.A0(\B_int[13] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][14] ), 
          .D1(GND_net), .CIN(n62303), .COUT(n62304), .S0(\m_cablesIn[18][14] ), 
          .S1(\m_cablesIn[18][15] ));
    defparam add_3537_15.INIT0 = 16'h6969;
    defparam add_3537_15.INIT1 = 16'h6969;
    defparam add_3537_15.INJECT1_0 = "NO";
    defparam add_3537_15.INJECT1_1 = "NO";
    CCU2D add_3537_13 (.A0(\B_int[11] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][12] ), 
          .D1(GND_net), .CIN(n62302), .COUT(n62303), .S0(\m_cablesIn[18][12] ), 
          .S1(\m_cablesIn[18][13] ));
    defparam add_3537_13.INIT0 = 16'h6969;
    defparam add_3537_13.INIT1 = 16'h6969;
    defparam add_3537_13.INJECT1_0 = "NO";
    defparam add_3537_13.INJECT1_1 = "NO";
    CCU2D add_3537_11 (.A0(\B_int[9] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][10] ), 
          .D1(GND_net), .CIN(n62301), .COUT(n62302), .S0(\m_cablesIn[18][10] ), 
          .S1(\m_cablesIn[18][11] ));
    defparam add_3537_11.INIT0 = 16'h6969;
    defparam add_3537_11.INIT1 = 16'h6969;
    defparam add_3537_11.INJECT1_0 = "NO";
    defparam add_3537_11.INJECT1_1 = "NO";
    CCU2D add_3537_9 (.A0(\B_int[7] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][8] ), 
          .D1(GND_net), .CIN(n62300), .COUT(n62301), .S0(\m_cablesIn[18][8] ), 
          .S1(\m_cablesIn[18][9] ));
    defparam add_3537_9.INIT0 = 16'h6969;
    defparam add_3537_9.INIT1 = 16'h6969;
    defparam add_3537_9.INJECT1_0 = "NO";
    defparam add_3537_9.INJECT1_1 = "NO";
    CCU2D add_3537_7 (.A0(\B_int[5] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][6] ), 
          .D1(GND_net), .CIN(n62299), .COUT(n62300), .S0(\m_cablesIn[18][6] ), 
          .S1(\m_cablesIn[18][7] ));
    defparam add_3537_7.INIT0 = 16'h6969;
    defparam add_3537_7.INIT1 = 16'h6969;
    defparam add_3537_7.INJECT1_0 = "NO";
    defparam add_3537_7.INJECT1_1 = "NO";
    CCU2D add_3537_5 (.A0(\B_int[3] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][4] ), 
          .D1(GND_net), .CIN(n62298), .COUT(n62299), .S0(\m_cablesIn[18][4] ), 
          .S1(\m_cablesIn[18][5] ));
    defparam add_3537_5.INIT0 = 16'h6969;
    defparam add_3537_5.INIT1 = 16'h6969;
    defparam add_3537_5.INJECT1_0 = "NO";
    defparam add_3537_5.INJECT1_1 = "NO";
    CCU2D add_3537_3 (.A0(\B_int[1] ), .B0(\QQ_in[17][16] ), .C0(\m_cablesIn[17][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[17][16] ), .C1(\m_cablesIn[17][2] ), 
          .D1(GND_net), .CIN(n62297), .COUT(n62298), .S0(\m_cablesIn[18][2] ), 
          .S1(\m_cablesIn[18][3] ));
    defparam add_3537_3.INIT0 = 16'h6969;
    defparam add_3537_3.INIT1 = 16'h6969;
    defparam add_3537_3.INJECT1_0 = "NO";
    defparam add_3537_3.INJECT1_1 = "NO";
    CCU2D add_3537_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[17][16] ), .C1(\frac_div[10] ), 
          .D1(GND_net), .COUT(n62297), .S1(\m_cablesIn[18][1] ));
    defparam add_3537_1.INIT0 = 16'hF000;
    defparam add_3537_1.INIT1 = 16'h6969;
    defparam add_3537_1.INJECT1_0 = "NO";
    defparam add_3537_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U17 
//

module \a_s(24)_U17  (\m_cablesIn[16][23] , \QQ_in[16][15] , GND_net, 
            \m_cablesIn[16][24] , \m_cablesIn[17][24] , \QQ_in[17][16] , 
            \B_int[21] , \m_cablesIn[16][21] , \B_int[22] , \m_cablesIn[16][22] , 
            \m_cablesIn[17][22] , \m_cablesIn[17][23] , \B_int[19] , \m_cablesIn[16][19] , 
            \B_int[20] , \m_cablesIn[16][20] , \m_cablesIn[17][20] , \m_cablesIn[17][21] , 
            \B_int[17] , \m_cablesIn[16][17] , \B_int[18] , \m_cablesIn[16][18] , 
            \m_cablesIn[17][18] , \m_cablesIn[17][19] , \B_int[15] , \m_cablesIn[16][15] , 
            \B_int[16] , \m_cablesIn[16][16] , \m_cablesIn[17][16] , \m_cablesIn[17][17] , 
            \B_int[13] , \m_cablesIn[16][13] , \B_int[14] , \m_cablesIn[16][14] , 
            \m_cablesIn[17][14] , \m_cablesIn[17][15] , \B_int[11] , \m_cablesIn[16][11] , 
            \B_int[12] , \m_cablesIn[16][12] , \m_cablesIn[17][12] , \m_cablesIn[17][13] , 
            \B_int[9] , \m_cablesIn[16][9] , \B_int[10] , \m_cablesIn[16][10] , 
            \m_cablesIn[17][10] , \m_cablesIn[17][11] , \B_int[7] , \m_cablesIn[16][7] , 
            \B_int[8] , \m_cablesIn[16][8] , \m_cablesIn[17][8] , \m_cablesIn[17][9] , 
            \B_int[5] , \m_cablesIn[16][5] , \B_int[6] , \m_cablesIn[16][6] , 
            \m_cablesIn[17][6] , \m_cablesIn[17][7] , \B_int[3] , \m_cablesIn[16][3] , 
            \B_int[4] , \m_cablesIn[16][4] , \m_cablesIn[17][4] , \m_cablesIn[17][5] , 
            \B_int[1] , \m_cablesIn[16][1] , \B_int[2] , \m_cablesIn[16][2] , 
            \m_cablesIn[17][2] , \m_cablesIn[17][3] , \B_int[0] , \frac_div[11] , 
            \m_cablesIn[17][1] );
    input \m_cablesIn[16][23] ;
    input \QQ_in[16][15] ;
    input GND_net;
    input \m_cablesIn[16][24] ;
    output \m_cablesIn[17][24] ;
    output \QQ_in[17][16] ;
    input \B_int[21] ;
    input \m_cablesIn[16][21] ;
    input \B_int[22] ;
    input \m_cablesIn[16][22] ;
    output \m_cablesIn[17][22] ;
    output \m_cablesIn[17][23] ;
    input \B_int[19] ;
    input \m_cablesIn[16][19] ;
    input \B_int[20] ;
    input \m_cablesIn[16][20] ;
    output \m_cablesIn[17][20] ;
    output \m_cablesIn[17][21] ;
    input \B_int[17] ;
    input \m_cablesIn[16][17] ;
    input \B_int[18] ;
    input \m_cablesIn[16][18] ;
    output \m_cablesIn[17][18] ;
    output \m_cablesIn[17][19] ;
    input \B_int[15] ;
    input \m_cablesIn[16][15] ;
    input \B_int[16] ;
    input \m_cablesIn[16][16] ;
    output \m_cablesIn[17][16] ;
    output \m_cablesIn[17][17] ;
    input \B_int[13] ;
    input \m_cablesIn[16][13] ;
    input \B_int[14] ;
    input \m_cablesIn[16][14] ;
    output \m_cablesIn[17][14] ;
    output \m_cablesIn[17][15] ;
    input \B_int[11] ;
    input \m_cablesIn[16][11] ;
    input \B_int[12] ;
    input \m_cablesIn[16][12] ;
    output \m_cablesIn[17][12] ;
    output \m_cablesIn[17][13] ;
    input \B_int[9] ;
    input \m_cablesIn[16][9] ;
    input \B_int[10] ;
    input \m_cablesIn[16][10] ;
    output \m_cablesIn[17][10] ;
    output \m_cablesIn[17][11] ;
    input \B_int[7] ;
    input \m_cablesIn[16][7] ;
    input \B_int[8] ;
    input \m_cablesIn[16][8] ;
    output \m_cablesIn[17][8] ;
    output \m_cablesIn[17][9] ;
    input \B_int[5] ;
    input \m_cablesIn[16][5] ;
    input \B_int[6] ;
    input \m_cablesIn[16][6] ;
    output \m_cablesIn[17][6] ;
    output \m_cablesIn[17][7] ;
    input \B_int[3] ;
    input \m_cablesIn[16][3] ;
    input \B_int[4] ;
    input \m_cablesIn[16][4] ;
    output \m_cablesIn[17][4] ;
    output \m_cablesIn[17][5] ;
    input \B_int[1] ;
    input \m_cablesIn[16][1] ;
    input \B_int[2] ;
    input \m_cablesIn[16][2] ;
    output \m_cablesIn[17][2] ;
    output \m_cablesIn[17][3] ;
    input \B_int[0] ;
    input \frac_div[11] ;
    output \m_cablesIn[17][1] ;
    
    
    wire n62321, n62320, n62319, n62318, n62317, n62316, n62315, 
        n62314, n62313, n62312, n62311, n62310;
    
    CCU2D add_3511_25 (.A0(\m_cablesIn[16][23] ), .B0(\QQ_in[16][15] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[16][24] ), .B1(\QQ_in[16][15] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62321), .S0(\m_cablesIn[17][24] ), 
          .S1(\QQ_in[17][16] ));
    defparam add_3511_25.INIT0 = 16'h5666;
    defparam add_3511_25.INIT1 = 16'h5999;
    defparam add_3511_25.INJECT1_0 = "NO";
    defparam add_3511_25.INJECT1_1 = "NO";
    CCU2D add_3511_23 (.A0(\B_int[21] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][22] ), 
          .D1(GND_net), .CIN(n62320), .COUT(n62321), .S0(\m_cablesIn[17][22] ), 
          .S1(\m_cablesIn[17][23] ));
    defparam add_3511_23.INIT0 = 16'h6969;
    defparam add_3511_23.INIT1 = 16'h6969;
    defparam add_3511_23.INJECT1_0 = "NO";
    defparam add_3511_23.INJECT1_1 = "NO";
    CCU2D add_3511_21 (.A0(\B_int[19] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][20] ), 
          .D1(GND_net), .CIN(n62319), .COUT(n62320), .S0(\m_cablesIn[17][20] ), 
          .S1(\m_cablesIn[17][21] ));
    defparam add_3511_21.INIT0 = 16'h6969;
    defparam add_3511_21.INIT1 = 16'h6969;
    defparam add_3511_21.INJECT1_0 = "NO";
    defparam add_3511_21.INJECT1_1 = "NO";
    CCU2D add_3511_19 (.A0(\B_int[17] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][18] ), 
          .D1(GND_net), .CIN(n62318), .COUT(n62319), .S0(\m_cablesIn[17][18] ), 
          .S1(\m_cablesIn[17][19] ));
    defparam add_3511_19.INIT0 = 16'h6969;
    defparam add_3511_19.INIT1 = 16'h6969;
    defparam add_3511_19.INJECT1_0 = "NO";
    defparam add_3511_19.INJECT1_1 = "NO";
    CCU2D add_3511_17 (.A0(\B_int[15] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][16] ), 
          .D1(GND_net), .CIN(n62317), .COUT(n62318), .S0(\m_cablesIn[17][16] ), 
          .S1(\m_cablesIn[17][17] ));
    defparam add_3511_17.INIT0 = 16'h6969;
    defparam add_3511_17.INIT1 = 16'h6969;
    defparam add_3511_17.INJECT1_0 = "NO";
    defparam add_3511_17.INJECT1_1 = "NO";
    CCU2D add_3511_15 (.A0(\B_int[13] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][14] ), 
          .D1(GND_net), .CIN(n62316), .COUT(n62317), .S0(\m_cablesIn[17][14] ), 
          .S1(\m_cablesIn[17][15] ));
    defparam add_3511_15.INIT0 = 16'h6969;
    defparam add_3511_15.INIT1 = 16'h6969;
    defparam add_3511_15.INJECT1_0 = "NO";
    defparam add_3511_15.INJECT1_1 = "NO";
    CCU2D add_3511_13 (.A0(\B_int[11] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][12] ), 
          .D1(GND_net), .CIN(n62315), .COUT(n62316), .S0(\m_cablesIn[17][12] ), 
          .S1(\m_cablesIn[17][13] ));
    defparam add_3511_13.INIT0 = 16'h6969;
    defparam add_3511_13.INIT1 = 16'h6969;
    defparam add_3511_13.INJECT1_0 = "NO";
    defparam add_3511_13.INJECT1_1 = "NO";
    CCU2D add_3511_11 (.A0(\B_int[9] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][10] ), 
          .D1(GND_net), .CIN(n62314), .COUT(n62315), .S0(\m_cablesIn[17][10] ), 
          .S1(\m_cablesIn[17][11] ));
    defparam add_3511_11.INIT0 = 16'h6969;
    defparam add_3511_11.INIT1 = 16'h6969;
    defparam add_3511_11.INJECT1_0 = "NO";
    defparam add_3511_11.INJECT1_1 = "NO";
    CCU2D add_3511_9 (.A0(\B_int[7] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][8] ), 
          .D1(GND_net), .CIN(n62313), .COUT(n62314), .S0(\m_cablesIn[17][8] ), 
          .S1(\m_cablesIn[17][9] ));
    defparam add_3511_9.INIT0 = 16'h6969;
    defparam add_3511_9.INIT1 = 16'h6969;
    defparam add_3511_9.INJECT1_0 = "NO";
    defparam add_3511_9.INJECT1_1 = "NO";
    CCU2D add_3511_7 (.A0(\B_int[5] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][6] ), 
          .D1(GND_net), .CIN(n62312), .COUT(n62313), .S0(\m_cablesIn[17][6] ), 
          .S1(\m_cablesIn[17][7] ));
    defparam add_3511_7.INIT0 = 16'h6969;
    defparam add_3511_7.INIT1 = 16'h6969;
    defparam add_3511_7.INJECT1_0 = "NO";
    defparam add_3511_7.INJECT1_1 = "NO";
    CCU2D add_3511_5 (.A0(\B_int[3] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][4] ), 
          .D1(GND_net), .CIN(n62311), .COUT(n62312), .S0(\m_cablesIn[17][4] ), 
          .S1(\m_cablesIn[17][5] ));
    defparam add_3511_5.INIT0 = 16'h6969;
    defparam add_3511_5.INIT1 = 16'h6969;
    defparam add_3511_5.INJECT1_0 = "NO";
    defparam add_3511_5.INJECT1_1 = "NO";
    CCU2D add_3511_3 (.A0(\B_int[1] ), .B0(\QQ_in[16][15] ), .C0(\m_cablesIn[16][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[16][15] ), .C1(\m_cablesIn[16][2] ), 
          .D1(GND_net), .CIN(n62310), .COUT(n62311), .S0(\m_cablesIn[17][2] ), 
          .S1(\m_cablesIn[17][3] ));
    defparam add_3511_3.INIT0 = 16'h6969;
    defparam add_3511_3.INIT1 = 16'h6969;
    defparam add_3511_3.INJECT1_0 = "NO";
    defparam add_3511_3.INJECT1_1 = "NO";
    CCU2D add_3511_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[16][15] ), .C1(\frac_div[11] ), 
          .D1(GND_net), .COUT(n62310), .S1(\m_cablesIn[17][1] ));
    defparam add_3511_1.INIT0 = 16'hF000;
    defparam add_3511_1.INIT1 = 16'h6969;
    defparam add_3511_1.INJECT1_0 = "NO";
    defparam add_3511_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U18 
//

module \a_s(24)_U18  (\m_cablesIn[15][23] , \QQ_in[15][14] , GND_net, 
            \m_cablesIn[15][24] , \m_cablesIn[16][24] , \QQ_in[16][15] , 
            \B_int[21] , \m_cablesIn[15][21] , \B_int[22] , \m_cablesIn[15][22] , 
            \m_cablesIn[16][22] , \m_cablesIn[16][23] , \B_int[19] , \m_cablesIn[15][19] , 
            \B_int[20] , \m_cablesIn[15][20] , \m_cablesIn[16][20] , \m_cablesIn[16][21] , 
            \B_int[17] , \m_cablesIn[15][17] , \B_int[18] , \m_cablesIn[15][18] , 
            \m_cablesIn[16][18] , \m_cablesIn[16][19] , \B_int[15] , \m_cablesIn[15][15] , 
            \B_int[16] , \m_cablesIn[15][16] , \m_cablesIn[16][16] , \m_cablesIn[16][17] , 
            \B_int[13] , \m_cablesIn[15][13] , \B_int[14] , \m_cablesIn[15][14] , 
            \m_cablesIn[16][14] , \m_cablesIn[16][15] , \B_int[11] , \m_cablesIn[15][11] , 
            \B_int[12] , \m_cablesIn[15][12] , \m_cablesIn[16][12] , \m_cablesIn[16][13] , 
            \B_int[9] , \m_cablesIn[15][9] , \B_int[10] , \m_cablesIn[15][10] , 
            \m_cablesIn[16][10] , \m_cablesIn[16][11] , \B_int[7] , \m_cablesIn[15][7] , 
            \B_int[8] , \m_cablesIn[15][8] , \m_cablesIn[16][8] , \m_cablesIn[16][9] , 
            \B_int[5] , \m_cablesIn[15][5] , \B_int[6] , \m_cablesIn[15][6] , 
            \m_cablesIn[16][6] , \m_cablesIn[16][7] , \B_int[3] , \m_cablesIn[15][3] , 
            \B_int[4] , \m_cablesIn[15][4] , \m_cablesIn[16][4] , \m_cablesIn[16][5] , 
            \B_int[1] , \m_cablesIn[15][1] , \B_int[2] , \m_cablesIn[15][2] , 
            \m_cablesIn[16][2] , \m_cablesIn[16][3] , \B_int[0] , \frac_div[12] , 
            \m_cablesIn[16][1] );
    input \m_cablesIn[15][23] ;
    input \QQ_in[15][14] ;
    input GND_net;
    input \m_cablesIn[15][24] ;
    output \m_cablesIn[16][24] ;
    output \QQ_in[16][15] ;
    input \B_int[21] ;
    input \m_cablesIn[15][21] ;
    input \B_int[22] ;
    input \m_cablesIn[15][22] ;
    output \m_cablesIn[16][22] ;
    output \m_cablesIn[16][23] ;
    input \B_int[19] ;
    input \m_cablesIn[15][19] ;
    input \B_int[20] ;
    input \m_cablesIn[15][20] ;
    output \m_cablesIn[16][20] ;
    output \m_cablesIn[16][21] ;
    input \B_int[17] ;
    input \m_cablesIn[15][17] ;
    input \B_int[18] ;
    input \m_cablesIn[15][18] ;
    output \m_cablesIn[16][18] ;
    output \m_cablesIn[16][19] ;
    input \B_int[15] ;
    input \m_cablesIn[15][15] ;
    input \B_int[16] ;
    input \m_cablesIn[15][16] ;
    output \m_cablesIn[16][16] ;
    output \m_cablesIn[16][17] ;
    input \B_int[13] ;
    input \m_cablesIn[15][13] ;
    input \B_int[14] ;
    input \m_cablesIn[15][14] ;
    output \m_cablesIn[16][14] ;
    output \m_cablesIn[16][15] ;
    input \B_int[11] ;
    input \m_cablesIn[15][11] ;
    input \B_int[12] ;
    input \m_cablesIn[15][12] ;
    output \m_cablesIn[16][12] ;
    output \m_cablesIn[16][13] ;
    input \B_int[9] ;
    input \m_cablesIn[15][9] ;
    input \B_int[10] ;
    input \m_cablesIn[15][10] ;
    output \m_cablesIn[16][10] ;
    output \m_cablesIn[16][11] ;
    input \B_int[7] ;
    input \m_cablesIn[15][7] ;
    input \B_int[8] ;
    input \m_cablesIn[15][8] ;
    output \m_cablesIn[16][8] ;
    output \m_cablesIn[16][9] ;
    input \B_int[5] ;
    input \m_cablesIn[15][5] ;
    input \B_int[6] ;
    input \m_cablesIn[15][6] ;
    output \m_cablesIn[16][6] ;
    output \m_cablesIn[16][7] ;
    input \B_int[3] ;
    input \m_cablesIn[15][3] ;
    input \B_int[4] ;
    input \m_cablesIn[15][4] ;
    output \m_cablesIn[16][4] ;
    output \m_cablesIn[16][5] ;
    input \B_int[1] ;
    input \m_cablesIn[15][1] ;
    input \B_int[2] ;
    input \m_cablesIn[15][2] ;
    output \m_cablesIn[16][2] ;
    output \m_cablesIn[16][3] ;
    input \B_int[0] ;
    input \frac_div[12] ;
    output \m_cablesIn[16][1] ;
    
    
    wire n62334, n62333, n62332, n62331, n62330, n62329, n62328, 
        n62327, n62326, n62325, n62324, n62323;
    
    CCU2D add_3485_25 (.A0(\m_cablesIn[15][23] ), .B0(\QQ_in[15][14] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[15][24] ), .B1(\QQ_in[15][14] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62334), .S0(\m_cablesIn[16][24] ), 
          .S1(\QQ_in[16][15] ));
    defparam add_3485_25.INIT0 = 16'h5666;
    defparam add_3485_25.INIT1 = 16'h5999;
    defparam add_3485_25.INJECT1_0 = "NO";
    defparam add_3485_25.INJECT1_1 = "NO";
    CCU2D add_3485_23 (.A0(\B_int[21] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][22] ), 
          .D1(GND_net), .CIN(n62333), .COUT(n62334), .S0(\m_cablesIn[16][22] ), 
          .S1(\m_cablesIn[16][23] ));
    defparam add_3485_23.INIT0 = 16'h6969;
    defparam add_3485_23.INIT1 = 16'h6969;
    defparam add_3485_23.INJECT1_0 = "NO";
    defparam add_3485_23.INJECT1_1 = "NO";
    CCU2D add_3485_21 (.A0(\B_int[19] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][20] ), 
          .D1(GND_net), .CIN(n62332), .COUT(n62333), .S0(\m_cablesIn[16][20] ), 
          .S1(\m_cablesIn[16][21] ));
    defparam add_3485_21.INIT0 = 16'h6969;
    defparam add_3485_21.INIT1 = 16'h6969;
    defparam add_3485_21.INJECT1_0 = "NO";
    defparam add_3485_21.INJECT1_1 = "NO";
    CCU2D add_3485_19 (.A0(\B_int[17] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][18] ), 
          .D1(GND_net), .CIN(n62331), .COUT(n62332), .S0(\m_cablesIn[16][18] ), 
          .S1(\m_cablesIn[16][19] ));
    defparam add_3485_19.INIT0 = 16'h6969;
    defparam add_3485_19.INIT1 = 16'h6969;
    defparam add_3485_19.INJECT1_0 = "NO";
    defparam add_3485_19.INJECT1_1 = "NO";
    CCU2D add_3485_17 (.A0(\B_int[15] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][16] ), 
          .D1(GND_net), .CIN(n62330), .COUT(n62331), .S0(\m_cablesIn[16][16] ), 
          .S1(\m_cablesIn[16][17] ));
    defparam add_3485_17.INIT0 = 16'h6969;
    defparam add_3485_17.INIT1 = 16'h6969;
    defparam add_3485_17.INJECT1_0 = "NO";
    defparam add_3485_17.INJECT1_1 = "NO";
    CCU2D add_3485_15 (.A0(\B_int[13] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][14] ), 
          .D1(GND_net), .CIN(n62329), .COUT(n62330), .S0(\m_cablesIn[16][14] ), 
          .S1(\m_cablesIn[16][15] ));
    defparam add_3485_15.INIT0 = 16'h6969;
    defparam add_3485_15.INIT1 = 16'h6969;
    defparam add_3485_15.INJECT1_0 = "NO";
    defparam add_3485_15.INJECT1_1 = "NO";
    CCU2D add_3485_13 (.A0(\B_int[11] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][12] ), 
          .D1(GND_net), .CIN(n62328), .COUT(n62329), .S0(\m_cablesIn[16][12] ), 
          .S1(\m_cablesIn[16][13] ));
    defparam add_3485_13.INIT0 = 16'h6969;
    defparam add_3485_13.INIT1 = 16'h6969;
    defparam add_3485_13.INJECT1_0 = "NO";
    defparam add_3485_13.INJECT1_1 = "NO";
    CCU2D add_3485_11 (.A0(\B_int[9] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][10] ), 
          .D1(GND_net), .CIN(n62327), .COUT(n62328), .S0(\m_cablesIn[16][10] ), 
          .S1(\m_cablesIn[16][11] ));
    defparam add_3485_11.INIT0 = 16'h6969;
    defparam add_3485_11.INIT1 = 16'h6969;
    defparam add_3485_11.INJECT1_0 = "NO";
    defparam add_3485_11.INJECT1_1 = "NO";
    CCU2D add_3485_9 (.A0(\B_int[7] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][8] ), 
          .D1(GND_net), .CIN(n62326), .COUT(n62327), .S0(\m_cablesIn[16][8] ), 
          .S1(\m_cablesIn[16][9] ));
    defparam add_3485_9.INIT0 = 16'h6969;
    defparam add_3485_9.INIT1 = 16'h6969;
    defparam add_3485_9.INJECT1_0 = "NO";
    defparam add_3485_9.INJECT1_1 = "NO";
    CCU2D add_3485_7 (.A0(\B_int[5] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][6] ), 
          .D1(GND_net), .CIN(n62325), .COUT(n62326), .S0(\m_cablesIn[16][6] ), 
          .S1(\m_cablesIn[16][7] ));
    defparam add_3485_7.INIT0 = 16'h6969;
    defparam add_3485_7.INIT1 = 16'h6969;
    defparam add_3485_7.INJECT1_0 = "NO";
    defparam add_3485_7.INJECT1_1 = "NO";
    CCU2D add_3485_5 (.A0(\B_int[3] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][4] ), 
          .D1(GND_net), .CIN(n62324), .COUT(n62325), .S0(\m_cablesIn[16][4] ), 
          .S1(\m_cablesIn[16][5] ));
    defparam add_3485_5.INIT0 = 16'h6969;
    defparam add_3485_5.INIT1 = 16'h6969;
    defparam add_3485_5.INJECT1_0 = "NO";
    defparam add_3485_5.INJECT1_1 = "NO";
    CCU2D add_3485_3 (.A0(\B_int[1] ), .B0(\QQ_in[15][14] ), .C0(\m_cablesIn[15][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[15][14] ), .C1(\m_cablesIn[15][2] ), 
          .D1(GND_net), .CIN(n62323), .COUT(n62324), .S0(\m_cablesIn[16][2] ), 
          .S1(\m_cablesIn[16][3] ));
    defparam add_3485_3.INIT0 = 16'h6969;
    defparam add_3485_3.INIT1 = 16'h6969;
    defparam add_3485_3.INJECT1_0 = "NO";
    defparam add_3485_3.INJECT1_1 = "NO";
    CCU2D add_3485_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[15][14] ), .C1(\frac_div[12] ), 
          .D1(GND_net), .COUT(n62323), .S1(\m_cablesIn[16][1] ));
    defparam add_3485_1.INIT0 = 16'hF000;
    defparam add_3485_1.INIT1 = 16'h6969;
    defparam add_3485_1.INJECT1_0 = "NO";
    defparam add_3485_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U19 
//

module \a_s(24)_U19  (\m_cablesIn[14][23] , \QQ_in[14][13] , GND_net, 
            \m_cablesIn[14][24] , \m_cablesIn[15][24] , \QQ_in[15][14] , 
            \B_int[21] , \m_cablesIn[14][21] , \B_int[22] , \m_cablesIn[14][22] , 
            \m_cablesIn[15][22] , \m_cablesIn[15][23] , \B_int[19] , \m_cablesIn[14][19] , 
            \B_int[20] , \m_cablesIn[14][20] , \m_cablesIn[15][20] , \m_cablesIn[15][21] , 
            \B_int[17] , \m_cablesIn[14][17] , \B_int[18] , \m_cablesIn[14][18] , 
            \m_cablesIn[15][18] , \m_cablesIn[15][19] , \B_int[15] , \m_cablesIn[14][15] , 
            \B_int[16] , \m_cablesIn[14][16] , \m_cablesIn[15][16] , \m_cablesIn[15][17] , 
            \B_int[13] , \m_cablesIn[14][13] , \B_int[14] , \m_cablesIn[14][14] , 
            \m_cablesIn[15][14] , \m_cablesIn[15][15] , \B_int[11] , \m_cablesIn[14][11] , 
            \B_int[12] , \m_cablesIn[14][12] , \m_cablesIn[15][12] , \m_cablesIn[15][13] , 
            \B_int[9] , \m_cablesIn[14][9] , \B_int[10] , \m_cablesIn[14][10] , 
            \m_cablesIn[15][10] , \m_cablesIn[15][11] , \B_int[7] , \m_cablesIn[14][7] , 
            \B_int[8] , \m_cablesIn[14][8] , \m_cablesIn[15][8] , \m_cablesIn[15][9] , 
            \B_int[5] , \m_cablesIn[14][5] , \B_int[6] , \m_cablesIn[14][6] , 
            \m_cablesIn[15][6] , \m_cablesIn[15][7] , \B_int[3] , \m_cablesIn[14][3] , 
            \B_int[4] , \m_cablesIn[14][4] , \m_cablesIn[15][4] , \m_cablesIn[15][5] , 
            \B_int[1] , \m_cablesIn[14][1] , \B_int[2] , \m_cablesIn[14][2] , 
            \m_cablesIn[15][2] , \m_cablesIn[15][3] , \B_int[0] , \frac_div[13] , 
            \m_cablesIn[15][1] );
    input \m_cablesIn[14][23] ;
    input \QQ_in[14][13] ;
    input GND_net;
    input \m_cablesIn[14][24] ;
    output \m_cablesIn[15][24] ;
    output \QQ_in[15][14] ;
    input \B_int[21] ;
    input \m_cablesIn[14][21] ;
    input \B_int[22] ;
    input \m_cablesIn[14][22] ;
    output \m_cablesIn[15][22] ;
    output \m_cablesIn[15][23] ;
    input \B_int[19] ;
    input \m_cablesIn[14][19] ;
    input \B_int[20] ;
    input \m_cablesIn[14][20] ;
    output \m_cablesIn[15][20] ;
    output \m_cablesIn[15][21] ;
    input \B_int[17] ;
    input \m_cablesIn[14][17] ;
    input \B_int[18] ;
    input \m_cablesIn[14][18] ;
    output \m_cablesIn[15][18] ;
    output \m_cablesIn[15][19] ;
    input \B_int[15] ;
    input \m_cablesIn[14][15] ;
    input \B_int[16] ;
    input \m_cablesIn[14][16] ;
    output \m_cablesIn[15][16] ;
    output \m_cablesIn[15][17] ;
    input \B_int[13] ;
    input \m_cablesIn[14][13] ;
    input \B_int[14] ;
    input \m_cablesIn[14][14] ;
    output \m_cablesIn[15][14] ;
    output \m_cablesIn[15][15] ;
    input \B_int[11] ;
    input \m_cablesIn[14][11] ;
    input \B_int[12] ;
    input \m_cablesIn[14][12] ;
    output \m_cablesIn[15][12] ;
    output \m_cablesIn[15][13] ;
    input \B_int[9] ;
    input \m_cablesIn[14][9] ;
    input \B_int[10] ;
    input \m_cablesIn[14][10] ;
    output \m_cablesIn[15][10] ;
    output \m_cablesIn[15][11] ;
    input \B_int[7] ;
    input \m_cablesIn[14][7] ;
    input \B_int[8] ;
    input \m_cablesIn[14][8] ;
    output \m_cablesIn[15][8] ;
    output \m_cablesIn[15][9] ;
    input \B_int[5] ;
    input \m_cablesIn[14][5] ;
    input \B_int[6] ;
    input \m_cablesIn[14][6] ;
    output \m_cablesIn[15][6] ;
    output \m_cablesIn[15][7] ;
    input \B_int[3] ;
    input \m_cablesIn[14][3] ;
    input \B_int[4] ;
    input \m_cablesIn[14][4] ;
    output \m_cablesIn[15][4] ;
    output \m_cablesIn[15][5] ;
    input \B_int[1] ;
    input \m_cablesIn[14][1] ;
    input \B_int[2] ;
    input \m_cablesIn[14][2] ;
    output \m_cablesIn[15][2] ;
    output \m_cablesIn[15][3] ;
    input \B_int[0] ;
    input \frac_div[13] ;
    output \m_cablesIn[15][1] ;
    
    
    wire n62347, n62346, n62345, n62344, n62343, n62342, n62341, 
        n62340, n62339, n62338, n62337, n62336;
    
    CCU2D add_3459_25 (.A0(\m_cablesIn[14][23] ), .B0(\QQ_in[14][13] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[14][24] ), .B1(\QQ_in[14][13] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62347), .S0(\m_cablesIn[15][24] ), 
          .S1(\QQ_in[15][14] ));
    defparam add_3459_25.INIT0 = 16'h5666;
    defparam add_3459_25.INIT1 = 16'h5999;
    defparam add_3459_25.INJECT1_0 = "NO";
    defparam add_3459_25.INJECT1_1 = "NO";
    CCU2D add_3459_23 (.A0(\B_int[21] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][22] ), 
          .D1(GND_net), .CIN(n62346), .COUT(n62347), .S0(\m_cablesIn[15][22] ), 
          .S1(\m_cablesIn[15][23] ));
    defparam add_3459_23.INIT0 = 16'h6969;
    defparam add_3459_23.INIT1 = 16'h6969;
    defparam add_3459_23.INJECT1_0 = "NO";
    defparam add_3459_23.INJECT1_1 = "NO";
    CCU2D add_3459_21 (.A0(\B_int[19] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][20] ), 
          .D1(GND_net), .CIN(n62345), .COUT(n62346), .S0(\m_cablesIn[15][20] ), 
          .S1(\m_cablesIn[15][21] ));
    defparam add_3459_21.INIT0 = 16'h6969;
    defparam add_3459_21.INIT1 = 16'h6969;
    defparam add_3459_21.INJECT1_0 = "NO";
    defparam add_3459_21.INJECT1_1 = "NO";
    CCU2D add_3459_19 (.A0(\B_int[17] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][18] ), 
          .D1(GND_net), .CIN(n62344), .COUT(n62345), .S0(\m_cablesIn[15][18] ), 
          .S1(\m_cablesIn[15][19] ));
    defparam add_3459_19.INIT0 = 16'h6969;
    defparam add_3459_19.INIT1 = 16'h6969;
    defparam add_3459_19.INJECT1_0 = "NO";
    defparam add_3459_19.INJECT1_1 = "NO";
    CCU2D add_3459_17 (.A0(\B_int[15] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][16] ), 
          .D1(GND_net), .CIN(n62343), .COUT(n62344), .S0(\m_cablesIn[15][16] ), 
          .S1(\m_cablesIn[15][17] ));
    defparam add_3459_17.INIT0 = 16'h6969;
    defparam add_3459_17.INIT1 = 16'h6969;
    defparam add_3459_17.INJECT1_0 = "NO";
    defparam add_3459_17.INJECT1_1 = "NO";
    CCU2D add_3459_15 (.A0(\B_int[13] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][14] ), 
          .D1(GND_net), .CIN(n62342), .COUT(n62343), .S0(\m_cablesIn[15][14] ), 
          .S1(\m_cablesIn[15][15] ));
    defparam add_3459_15.INIT0 = 16'h6969;
    defparam add_3459_15.INIT1 = 16'h6969;
    defparam add_3459_15.INJECT1_0 = "NO";
    defparam add_3459_15.INJECT1_1 = "NO";
    CCU2D add_3459_13 (.A0(\B_int[11] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][12] ), 
          .D1(GND_net), .CIN(n62341), .COUT(n62342), .S0(\m_cablesIn[15][12] ), 
          .S1(\m_cablesIn[15][13] ));
    defparam add_3459_13.INIT0 = 16'h6969;
    defparam add_3459_13.INIT1 = 16'h6969;
    defparam add_3459_13.INJECT1_0 = "NO";
    defparam add_3459_13.INJECT1_1 = "NO";
    CCU2D add_3459_11 (.A0(\B_int[9] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][10] ), 
          .D1(GND_net), .CIN(n62340), .COUT(n62341), .S0(\m_cablesIn[15][10] ), 
          .S1(\m_cablesIn[15][11] ));
    defparam add_3459_11.INIT0 = 16'h6969;
    defparam add_3459_11.INIT1 = 16'h6969;
    defparam add_3459_11.INJECT1_0 = "NO";
    defparam add_3459_11.INJECT1_1 = "NO";
    CCU2D add_3459_9 (.A0(\B_int[7] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][8] ), 
          .D1(GND_net), .CIN(n62339), .COUT(n62340), .S0(\m_cablesIn[15][8] ), 
          .S1(\m_cablesIn[15][9] ));
    defparam add_3459_9.INIT0 = 16'h6969;
    defparam add_3459_9.INIT1 = 16'h6969;
    defparam add_3459_9.INJECT1_0 = "NO";
    defparam add_3459_9.INJECT1_1 = "NO";
    CCU2D add_3459_7 (.A0(\B_int[5] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][6] ), 
          .D1(GND_net), .CIN(n62338), .COUT(n62339), .S0(\m_cablesIn[15][6] ), 
          .S1(\m_cablesIn[15][7] ));
    defparam add_3459_7.INIT0 = 16'h6969;
    defparam add_3459_7.INIT1 = 16'h6969;
    defparam add_3459_7.INJECT1_0 = "NO";
    defparam add_3459_7.INJECT1_1 = "NO";
    CCU2D add_3459_5 (.A0(\B_int[3] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][4] ), 
          .D1(GND_net), .CIN(n62337), .COUT(n62338), .S0(\m_cablesIn[15][4] ), 
          .S1(\m_cablesIn[15][5] ));
    defparam add_3459_5.INIT0 = 16'h6969;
    defparam add_3459_5.INIT1 = 16'h6969;
    defparam add_3459_5.INJECT1_0 = "NO";
    defparam add_3459_5.INJECT1_1 = "NO";
    CCU2D add_3459_3 (.A0(\B_int[1] ), .B0(\QQ_in[14][13] ), .C0(\m_cablesIn[14][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[14][13] ), .C1(\m_cablesIn[14][2] ), 
          .D1(GND_net), .CIN(n62336), .COUT(n62337), .S0(\m_cablesIn[15][2] ), 
          .S1(\m_cablesIn[15][3] ));
    defparam add_3459_3.INIT0 = 16'h6969;
    defparam add_3459_3.INIT1 = 16'h6969;
    defparam add_3459_3.INJECT1_0 = "NO";
    defparam add_3459_3.INJECT1_1 = "NO";
    CCU2D add_3459_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[14][13] ), .C1(\frac_div[13] ), 
          .D1(GND_net), .COUT(n62336), .S1(\m_cablesIn[15][1] ));
    defparam add_3459_1.INIT0 = 16'hF000;
    defparam add_3459_1.INIT1 = 16'h6969;
    defparam add_3459_1.INJECT1_0 = "NO";
    defparam add_3459_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U20 
//

module \a_s(24)_U20  (\m_cablesIn[13][23] , \QQ_in[13][12] , GND_net, 
            \m_cablesIn[13][24] , \m_cablesIn[14][24] , \QQ_in[14][13] , 
            \B_int[21] , \m_cablesIn[13][21] , \B_int[22] , \m_cablesIn[13][22] , 
            \m_cablesIn[14][22] , \m_cablesIn[14][23] , \B_int[19] , \m_cablesIn[13][19] , 
            \B_int[20] , \m_cablesIn[13][20] , \m_cablesIn[14][20] , \m_cablesIn[14][21] , 
            \B_int[17] , \m_cablesIn[13][17] , \B_int[18] , \m_cablesIn[13][18] , 
            \m_cablesIn[14][18] , \m_cablesIn[14][19] , \B_int[15] , \m_cablesIn[13][15] , 
            \B_int[16] , \m_cablesIn[13][16] , \m_cablesIn[14][16] , \m_cablesIn[14][17] , 
            \B_int[13] , \m_cablesIn[13][13] , \B_int[14] , \m_cablesIn[13][14] , 
            \m_cablesIn[14][14] , \m_cablesIn[14][15] , \B_int[11] , \m_cablesIn[13][11] , 
            \B_int[12] , \m_cablesIn[13][12] , \m_cablesIn[14][12] , \m_cablesIn[14][13] , 
            \B_int[9] , \m_cablesIn[13][9] , \B_int[10] , \m_cablesIn[13][10] , 
            \m_cablesIn[14][10] , \m_cablesIn[14][11] , \B_int[7] , \m_cablesIn[13][7] , 
            \B_int[8] , \m_cablesIn[13][8] , \m_cablesIn[14][8] , \m_cablesIn[14][9] , 
            \B_int[5] , \m_cablesIn[13][5] , \B_int[6] , \m_cablesIn[13][6] , 
            \m_cablesIn[14][6] , \m_cablesIn[14][7] , \B_int[3] , \m_cablesIn[13][3] , 
            \B_int[4] , \m_cablesIn[13][4] , \m_cablesIn[14][4] , \m_cablesIn[14][5] , 
            \B_int[1] , \m_cablesIn[13][1] , \B_int[2] , \m_cablesIn[13][2] , 
            \m_cablesIn[14][2] , \m_cablesIn[14][3] , \B_int[0] , \frac_div[14] , 
            \m_cablesIn[14][1] );
    input \m_cablesIn[13][23] ;
    input \QQ_in[13][12] ;
    input GND_net;
    input \m_cablesIn[13][24] ;
    output \m_cablesIn[14][24] ;
    output \QQ_in[14][13] ;
    input \B_int[21] ;
    input \m_cablesIn[13][21] ;
    input \B_int[22] ;
    input \m_cablesIn[13][22] ;
    output \m_cablesIn[14][22] ;
    output \m_cablesIn[14][23] ;
    input \B_int[19] ;
    input \m_cablesIn[13][19] ;
    input \B_int[20] ;
    input \m_cablesIn[13][20] ;
    output \m_cablesIn[14][20] ;
    output \m_cablesIn[14][21] ;
    input \B_int[17] ;
    input \m_cablesIn[13][17] ;
    input \B_int[18] ;
    input \m_cablesIn[13][18] ;
    output \m_cablesIn[14][18] ;
    output \m_cablesIn[14][19] ;
    input \B_int[15] ;
    input \m_cablesIn[13][15] ;
    input \B_int[16] ;
    input \m_cablesIn[13][16] ;
    output \m_cablesIn[14][16] ;
    output \m_cablesIn[14][17] ;
    input \B_int[13] ;
    input \m_cablesIn[13][13] ;
    input \B_int[14] ;
    input \m_cablesIn[13][14] ;
    output \m_cablesIn[14][14] ;
    output \m_cablesIn[14][15] ;
    input \B_int[11] ;
    input \m_cablesIn[13][11] ;
    input \B_int[12] ;
    input \m_cablesIn[13][12] ;
    output \m_cablesIn[14][12] ;
    output \m_cablesIn[14][13] ;
    input \B_int[9] ;
    input \m_cablesIn[13][9] ;
    input \B_int[10] ;
    input \m_cablesIn[13][10] ;
    output \m_cablesIn[14][10] ;
    output \m_cablesIn[14][11] ;
    input \B_int[7] ;
    input \m_cablesIn[13][7] ;
    input \B_int[8] ;
    input \m_cablesIn[13][8] ;
    output \m_cablesIn[14][8] ;
    output \m_cablesIn[14][9] ;
    input \B_int[5] ;
    input \m_cablesIn[13][5] ;
    input \B_int[6] ;
    input \m_cablesIn[13][6] ;
    output \m_cablesIn[14][6] ;
    output \m_cablesIn[14][7] ;
    input \B_int[3] ;
    input \m_cablesIn[13][3] ;
    input \B_int[4] ;
    input \m_cablesIn[13][4] ;
    output \m_cablesIn[14][4] ;
    output \m_cablesIn[14][5] ;
    input \B_int[1] ;
    input \m_cablesIn[13][1] ;
    input \B_int[2] ;
    input \m_cablesIn[13][2] ;
    output \m_cablesIn[14][2] ;
    output \m_cablesIn[14][3] ;
    input \B_int[0] ;
    input \frac_div[14] ;
    output \m_cablesIn[14][1] ;
    
    
    wire n62360, n62359, n62358, n62357, n62356, n62355, n62354, 
        n62353, n62352, n62351, n62350, n62349;
    
    CCU2D add_3433_25 (.A0(\m_cablesIn[13][23] ), .B0(\QQ_in[13][12] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[13][24] ), .B1(\QQ_in[13][12] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62360), .S0(\m_cablesIn[14][24] ), 
          .S1(\QQ_in[14][13] ));
    defparam add_3433_25.INIT0 = 16'h5666;
    defparam add_3433_25.INIT1 = 16'h5999;
    defparam add_3433_25.INJECT1_0 = "NO";
    defparam add_3433_25.INJECT1_1 = "NO";
    CCU2D add_3433_23 (.A0(\B_int[21] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][22] ), 
          .D1(GND_net), .CIN(n62359), .COUT(n62360), .S0(\m_cablesIn[14][22] ), 
          .S1(\m_cablesIn[14][23] ));
    defparam add_3433_23.INIT0 = 16'h6969;
    defparam add_3433_23.INIT1 = 16'h6969;
    defparam add_3433_23.INJECT1_0 = "NO";
    defparam add_3433_23.INJECT1_1 = "NO";
    CCU2D add_3433_21 (.A0(\B_int[19] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][20] ), 
          .D1(GND_net), .CIN(n62358), .COUT(n62359), .S0(\m_cablesIn[14][20] ), 
          .S1(\m_cablesIn[14][21] ));
    defparam add_3433_21.INIT0 = 16'h6969;
    defparam add_3433_21.INIT1 = 16'h6969;
    defparam add_3433_21.INJECT1_0 = "NO";
    defparam add_3433_21.INJECT1_1 = "NO";
    CCU2D add_3433_19 (.A0(\B_int[17] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][18] ), 
          .D1(GND_net), .CIN(n62357), .COUT(n62358), .S0(\m_cablesIn[14][18] ), 
          .S1(\m_cablesIn[14][19] ));
    defparam add_3433_19.INIT0 = 16'h6969;
    defparam add_3433_19.INIT1 = 16'h6969;
    defparam add_3433_19.INJECT1_0 = "NO";
    defparam add_3433_19.INJECT1_1 = "NO";
    CCU2D add_3433_17 (.A0(\B_int[15] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][16] ), 
          .D1(GND_net), .CIN(n62356), .COUT(n62357), .S0(\m_cablesIn[14][16] ), 
          .S1(\m_cablesIn[14][17] ));
    defparam add_3433_17.INIT0 = 16'h6969;
    defparam add_3433_17.INIT1 = 16'h6969;
    defparam add_3433_17.INJECT1_0 = "NO";
    defparam add_3433_17.INJECT1_1 = "NO";
    CCU2D add_3433_15 (.A0(\B_int[13] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][14] ), 
          .D1(GND_net), .CIN(n62355), .COUT(n62356), .S0(\m_cablesIn[14][14] ), 
          .S1(\m_cablesIn[14][15] ));
    defparam add_3433_15.INIT0 = 16'h6969;
    defparam add_3433_15.INIT1 = 16'h6969;
    defparam add_3433_15.INJECT1_0 = "NO";
    defparam add_3433_15.INJECT1_1 = "NO";
    CCU2D add_3433_13 (.A0(\B_int[11] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][12] ), 
          .D1(GND_net), .CIN(n62354), .COUT(n62355), .S0(\m_cablesIn[14][12] ), 
          .S1(\m_cablesIn[14][13] ));
    defparam add_3433_13.INIT0 = 16'h6969;
    defparam add_3433_13.INIT1 = 16'h6969;
    defparam add_3433_13.INJECT1_0 = "NO";
    defparam add_3433_13.INJECT1_1 = "NO";
    CCU2D add_3433_11 (.A0(\B_int[9] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][10] ), 
          .D1(GND_net), .CIN(n62353), .COUT(n62354), .S0(\m_cablesIn[14][10] ), 
          .S1(\m_cablesIn[14][11] ));
    defparam add_3433_11.INIT0 = 16'h6969;
    defparam add_3433_11.INIT1 = 16'h6969;
    defparam add_3433_11.INJECT1_0 = "NO";
    defparam add_3433_11.INJECT1_1 = "NO";
    CCU2D add_3433_9 (.A0(\B_int[7] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][8] ), 
          .D1(GND_net), .CIN(n62352), .COUT(n62353), .S0(\m_cablesIn[14][8] ), 
          .S1(\m_cablesIn[14][9] ));
    defparam add_3433_9.INIT0 = 16'h6969;
    defparam add_3433_9.INIT1 = 16'h6969;
    defparam add_3433_9.INJECT1_0 = "NO";
    defparam add_3433_9.INJECT1_1 = "NO";
    CCU2D add_3433_7 (.A0(\B_int[5] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][6] ), 
          .D1(GND_net), .CIN(n62351), .COUT(n62352), .S0(\m_cablesIn[14][6] ), 
          .S1(\m_cablesIn[14][7] ));
    defparam add_3433_7.INIT0 = 16'h6969;
    defparam add_3433_7.INIT1 = 16'h6969;
    defparam add_3433_7.INJECT1_0 = "NO";
    defparam add_3433_7.INJECT1_1 = "NO";
    CCU2D add_3433_5 (.A0(\B_int[3] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][4] ), 
          .D1(GND_net), .CIN(n62350), .COUT(n62351), .S0(\m_cablesIn[14][4] ), 
          .S1(\m_cablesIn[14][5] ));
    defparam add_3433_5.INIT0 = 16'h6969;
    defparam add_3433_5.INIT1 = 16'h6969;
    defparam add_3433_5.INJECT1_0 = "NO";
    defparam add_3433_5.INJECT1_1 = "NO";
    CCU2D add_3433_3 (.A0(\B_int[1] ), .B0(\QQ_in[13][12] ), .C0(\m_cablesIn[13][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[13][12] ), .C1(\m_cablesIn[13][2] ), 
          .D1(GND_net), .CIN(n62349), .COUT(n62350), .S0(\m_cablesIn[14][2] ), 
          .S1(\m_cablesIn[14][3] ));
    defparam add_3433_3.INIT0 = 16'h6969;
    defparam add_3433_3.INIT1 = 16'h6969;
    defparam add_3433_3.INJECT1_0 = "NO";
    defparam add_3433_3.INJECT1_1 = "NO";
    CCU2D add_3433_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[13][12] ), .C1(\frac_div[14] ), 
          .D1(GND_net), .COUT(n62349), .S1(\m_cablesIn[14][1] ));
    defparam add_3433_1.INIT0 = 16'hF000;
    defparam add_3433_1.INIT1 = 16'h6969;
    defparam add_3433_1.INJECT1_0 = "NO";
    defparam add_3433_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U21 
//

module \a_s(24)_U21  (\m_cablesIn[12][23] , \QQ_in[12][11] , GND_net, 
            \m_cablesIn[12][24] , \m_cablesIn[13][24] , \QQ_in[13][12] , 
            \B_int[21] , \m_cablesIn[12][21] , \B_int[22] , \m_cablesIn[12][22] , 
            \m_cablesIn[13][22] , \m_cablesIn[13][23] , \B_int[19] , \m_cablesIn[12][19] , 
            \B_int[20] , \m_cablesIn[12][20] , \m_cablesIn[13][20] , \m_cablesIn[13][21] , 
            \B_int[17] , \m_cablesIn[12][17] , \B_int[18] , \m_cablesIn[12][18] , 
            \m_cablesIn[13][18] , \m_cablesIn[13][19] , \B_int[15] , \m_cablesIn[12][15] , 
            \B_int[16] , \m_cablesIn[12][16] , \m_cablesIn[13][16] , \m_cablesIn[13][17] , 
            \B_int[13] , \m_cablesIn[12][13] , \B_int[14] , \m_cablesIn[12][14] , 
            \m_cablesIn[13][14] , \m_cablesIn[13][15] , \B_int[11] , \m_cablesIn[12][11] , 
            \B_int[12] , \m_cablesIn[12][12] , \m_cablesIn[13][12] , \m_cablesIn[13][13] , 
            \B_int[9] , \m_cablesIn[12][9] , \B_int[10] , \m_cablesIn[12][10] , 
            \m_cablesIn[13][10] , \m_cablesIn[13][11] , \B_int[7] , \m_cablesIn[12][7] , 
            \B_int[8] , \m_cablesIn[12][8] , \m_cablesIn[13][8] , \m_cablesIn[13][9] , 
            \B_int[5] , \m_cablesIn[12][5] , \B_int[6] , \m_cablesIn[12][6] , 
            \m_cablesIn[13][6] , \m_cablesIn[13][7] , \B_int[3] , \m_cablesIn[12][3] , 
            \B_int[4] , \m_cablesIn[12][4] , \m_cablesIn[13][4] , \m_cablesIn[13][5] , 
            \B_int[1] , \m_cablesIn[12][1] , \B_int[2] , \m_cablesIn[12][2] , 
            \m_cablesIn[13][2] , \m_cablesIn[13][3] , \B_int[0] , \frac_div[15] , 
            \m_cablesIn[13][1] );
    input \m_cablesIn[12][23] ;
    input \QQ_in[12][11] ;
    input GND_net;
    input \m_cablesIn[12][24] ;
    output \m_cablesIn[13][24] ;
    output \QQ_in[13][12] ;
    input \B_int[21] ;
    input \m_cablesIn[12][21] ;
    input \B_int[22] ;
    input \m_cablesIn[12][22] ;
    output \m_cablesIn[13][22] ;
    output \m_cablesIn[13][23] ;
    input \B_int[19] ;
    input \m_cablesIn[12][19] ;
    input \B_int[20] ;
    input \m_cablesIn[12][20] ;
    output \m_cablesIn[13][20] ;
    output \m_cablesIn[13][21] ;
    input \B_int[17] ;
    input \m_cablesIn[12][17] ;
    input \B_int[18] ;
    input \m_cablesIn[12][18] ;
    output \m_cablesIn[13][18] ;
    output \m_cablesIn[13][19] ;
    input \B_int[15] ;
    input \m_cablesIn[12][15] ;
    input \B_int[16] ;
    input \m_cablesIn[12][16] ;
    output \m_cablesIn[13][16] ;
    output \m_cablesIn[13][17] ;
    input \B_int[13] ;
    input \m_cablesIn[12][13] ;
    input \B_int[14] ;
    input \m_cablesIn[12][14] ;
    output \m_cablesIn[13][14] ;
    output \m_cablesIn[13][15] ;
    input \B_int[11] ;
    input \m_cablesIn[12][11] ;
    input \B_int[12] ;
    input \m_cablesIn[12][12] ;
    output \m_cablesIn[13][12] ;
    output \m_cablesIn[13][13] ;
    input \B_int[9] ;
    input \m_cablesIn[12][9] ;
    input \B_int[10] ;
    input \m_cablesIn[12][10] ;
    output \m_cablesIn[13][10] ;
    output \m_cablesIn[13][11] ;
    input \B_int[7] ;
    input \m_cablesIn[12][7] ;
    input \B_int[8] ;
    input \m_cablesIn[12][8] ;
    output \m_cablesIn[13][8] ;
    output \m_cablesIn[13][9] ;
    input \B_int[5] ;
    input \m_cablesIn[12][5] ;
    input \B_int[6] ;
    input \m_cablesIn[12][6] ;
    output \m_cablesIn[13][6] ;
    output \m_cablesIn[13][7] ;
    input \B_int[3] ;
    input \m_cablesIn[12][3] ;
    input \B_int[4] ;
    input \m_cablesIn[12][4] ;
    output \m_cablesIn[13][4] ;
    output \m_cablesIn[13][5] ;
    input \B_int[1] ;
    input \m_cablesIn[12][1] ;
    input \B_int[2] ;
    input \m_cablesIn[12][2] ;
    output \m_cablesIn[13][2] ;
    output \m_cablesIn[13][3] ;
    input \B_int[0] ;
    input \frac_div[15] ;
    output \m_cablesIn[13][1] ;
    
    
    wire n62373, n62372, n62371, n62370, n62369, n62368, n62367, 
        n62366, n62365, n62364, n62363, n62362;
    
    CCU2D add_3407_25 (.A0(\m_cablesIn[12][23] ), .B0(\QQ_in[12][11] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[12][24] ), .B1(\QQ_in[12][11] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62373), .S0(\m_cablesIn[13][24] ), 
          .S1(\QQ_in[13][12] ));
    defparam add_3407_25.INIT0 = 16'h5666;
    defparam add_3407_25.INIT1 = 16'h5999;
    defparam add_3407_25.INJECT1_0 = "NO";
    defparam add_3407_25.INJECT1_1 = "NO";
    CCU2D add_3407_23 (.A0(\B_int[21] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][22] ), 
          .D1(GND_net), .CIN(n62372), .COUT(n62373), .S0(\m_cablesIn[13][22] ), 
          .S1(\m_cablesIn[13][23] ));
    defparam add_3407_23.INIT0 = 16'h6969;
    defparam add_3407_23.INIT1 = 16'h6969;
    defparam add_3407_23.INJECT1_0 = "NO";
    defparam add_3407_23.INJECT1_1 = "NO";
    CCU2D add_3407_21 (.A0(\B_int[19] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][20] ), 
          .D1(GND_net), .CIN(n62371), .COUT(n62372), .S0(\m_cablesIn[13][20] ), 
          .S1(\m_cablesIn[13][21] ));
    defparam add_3407_21.INIT0 = 16'h6969;
    defparam add_3407_21.INIT1 = 16'h6969;
    defparam add_3407_21.INJECT1_0 = "NO";
    defparam add_3407_21.INJECT1_1 = "NO";
    CCU2D add_3407_19 (.A0(\B_int[17] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][18] ), 
          .D1(GND_net), .CIN(n62370), .COUT(n62371), .S0(\m_cablesIn[13][18] ), 
          .S1(\m_cablesIn[13][19] ));
    defparam add_3407_19.INIT0 = 16'h6969;
    defparam add_3407_19.INIT1 = 16'h6969;
    defparam add_3407_19.INJECT1_0 = "NO";
    defparam add_3407_19.INJECT1_1 = "NO";
    CCU2D add_3407_17 (.A0(\B_int[15] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][16] ), 
          .D1(GND_net), .CIN(n62369), .COUT(n62370), .S0(\m_cablesIn[13][16] ), 
          .S1(\m_cablesIn[13][17] ));
    defparam add_3407_17.INIT0 = 16'h6969;
    defparam add_3407_17.INIT1 = 16'h6969;
    defparam add_3407_17.INJECT1_0 = "NO";
    defparam add_3407_17.INJECT1_1 = "NO";
    CCU2D add_3407_15 (.A0(\B_int[13] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][14] ), 
          .D1(GND_net), .CIN(n62368), .COUT(n62369), .S0(\m_cablesIn[13][14] ), 
          .S1(\m_cablesIn[13][15] ));
    defparam add_3407_15.INIT0 = 16'h6969;
    defparam add_3407_15.INIT1 = 16'h6969;
    defparam add_3407_15.INJECT1_0 = "NO";
    defparam add_3407_15.INJECT1_1 = "NO";
    CCU2D add_3407_13 (.A0(\B_int[11] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][12] ), 
          .D1(GND_net), .CIN(n62367), .COUT(n62368), .S0(\m_cablesIn[13][12] ), 
          .S1(\m_cablesIn[13][13] ));
    defparam add_3407_13.INIT0 = 16'h6969;
    defparam add_3407_13.INIT1 = 16'h6969;
    defparam add_3407_13.INJECT1_0 = "NO";
    defparam add_3407_13.INJECT1_1 = "NO";
    CCU2D add_3407_11 (.A0(\B_int[9] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][10] ), 
          .D1(GND_net), .CIN(n62366), .COUT(n62367), .S0(\m_cablesIn[13][10] ), 
          .S1(\m_cablesIn[13][11] ));
    defparam add_3407_11.INIT0 = 16'h6969;
    defparam add_3407_11.INIT1 = 16'h6969;
    defparam add_3407_11.INJECT1_0 = "NO";
    defparam add_3407_11.INJECT1_1 = "NO";
    CCU2D add_3407_9 (.A0(\B_int[7] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][8] ), 
          .D1(GND_net), .CIN(n62365), .COUT(n62366), .S0(\m_cablesIn[13][8] ), 
          .S1(\m_cablesIn[13][9] ));
    defparam add_3407_9.INIT0 = 16'h6969;
    defparam add_3407_9.INIT1 = 16'h6969;
    defparam add_3407_9.INJECT1_0 = "NO";
    defparam add_3407_9.INJECT1_1 = "NO";
    CCU2D add_3407_7 (.A0(\B_int[5] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][6] ), 
          .D1(GND_net), .CIN(n62364), .COUT(n62365), .S0(\m_cablesIn[13][6] ), 
          .S1(\m_cablesIn[13][7] ));
    defparam add_3407_7.INIT0 = 16'h6969;
    defparam add_3407_7.INIT1 = 16'h6969;
    defparam add_3407_7.INJECT1_0 = "NO";
    defparam add_3407_7.INJECT1_1 = "NO";
    CCU2D add_3407_5 (.A0(\B_int[3] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][4] ), 
          .D1(GND_net), .CIN(n62363), .COUT(n62364), .S0(\m_cablesIn[13][4] ), 
          .S1(\m_cablesIn[13][5] ));
    defparam add_3407_5.INIT0 = 16'h6969;
    defparam add_3407_5.INIT1 = 16'h6969;
    defparam add_3407_5.INJECT1_0 = "NO";
    defparam add_3407_5.INJECT1_1 = "NO";
    CCU2D add_3407_3 (.A0(\B_int[1] ), .B0(\QQ_in[12][11] ), .C0(\m_cablesIn[12][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[12][11] ), .C1(\m_cablesIn[12][2] ), 
          .D1(GND_net), .CIN(n62362), .COUT(n62363), .S0(\m_cablesIn[13][2] ), 
          .S1(\m_cablesIn[13][3] ));
    defparam add_3407_3.INIT0 = 16'h6969;
    defparam add_3407_3.INIT1 = 16'h6969;
    defparam add_3407_3.INJECT1_0 = "NO";
    defparam add_3407_3.INJECT1_1 = "NO";
    CCU2D add_3407_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[12][11] ), .C1(\frac_div[15] ), 
          .D1(GND_net), .COUT(n62362), .S1(\m_cablesIn[13][1] ));
    defparam add_3407_1.INIT0 = 16'hF000;
    defparam add_3407_1.INIT1 = 16'h6969;
    defparam add_3407_1.INJECT1_0 = "NO";
    defparam add_3407_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U22 
//

module \a_s(24)_U22  (\m_cablesIn[11][23] , \QQ_in[11][10] , GND_net, 
            \m_cablesIn[11][24] , \m_cablesIn[12][24] , \QQ_in[12][11] , 
            \B_int[21] , \m_cablesIn[11][21] , \B_int[22] , \m_cablesIn[11][22] , 
            \m_cablesIn[12][22] , \m_cablesIn[12][23] , \B_int[19] , \m_cablesIn[11][19] , 
            \B_int[20] , \m_cablesIn[11][20] , \m_cablesIn[12][20] , \m_cablesIn[12][21] , 
            \B_int[17] , \m_cablesIn[11][17] , \B_int[18] , \m_cablesIn[11][18] , 
            \m_cablesIn[12][18] , \m_cablesIn[12][19] , \B_int[15] , \m_cablesIn[11][15] , 
            \B_int[16] , \m_cablesIn[11][16] , \m_cablesIn[12][16] , \m_cablesIn[12][17] , 
            \B_int[13] , \m_cablesIn[11][13] , \B_int[14] , \m_cablesIn[11][14] , 
            \m_cablesIn[12][14] , \m_cablesIn[12][15] , \B_int[11] , \m_cablesIn[11][11] , 
            \B_int[12] , \m_cablesIn[11][12] , \m_cablesIn[12][12] , \m_cablesIn[12][13] , 
            \B_int[9] , \m_cablesIn[11][9] , \B_int[10] , \m_cablesIn[11][10] , 
            \m_cablesIn[12][10] , \m_cablesIn[12][11] , \B_int[7] , \m_cablesIn[11][7] , 
            \B_int[8] , \m_cablesIn[11][8] , \m_cablesIn[12][8] , \m_cablesIn[12][9] , 
            \B_int[5] , \m_cablesIn[11][5] , \B_int[6] , \m_cablesIn[11][6] , 
            \m_cablesIn[12][6] , \m_cablesIn[12][7] , \B_int[3] , \m_cablesIn[11][3] , 
            \B_int[4] , \m_cablesIn[11][4] , \m_cablesIn[12][4] , \m_cablesIn[12][5] , 
            \B_int[1] , \m_cablesIn[11][1] , \B_int[2] , \m_cablesIn[11][2] , 
            \m_cablesIn[12][2] , \m_cablesIn[12][3] , \B_int[0] , \frac_div[16] , 
            \m_cablesIn[12][1] );
    input \m_cablesIn[11][23] ;
    input \QQ_in[11][10] ;
    input GND_net;
    input \m_cablesIn[11][24] ;
    output \m_cablesIn[12][24] ;
    output \QQ_in[12][11] ;
    input \B_int[21] ;
    input \m_cablesIn[11][21] ;
    input \B_int[22] ;
    input \m_cablesIn[11][22] ;
    output \m_cablesIn[12][22] ;
    output \m_cablesIn[12][23] ;
    input \B_int[19] ;
    input \m_cablesIn[11][19] ;
    input \B_int[20] ;
    input \m_cablesIn[11][20] ;
    output \m_cablesIn[12][20] ;
    output \m_cablesIn[12][21] ;
    input \B_int[17] ;
    input \m_cablesIn[11][17] ;
    input \B_int[18] ;
    input \m_cablesIn[11][18] ;
    output \m_cablesIn[12][18] ;
    output \m_cablesIn[12][19] ;
    input \B_int[15] ;
    input \m_cablesIn[11][15] ;
    input \B_int[16] ;
    input \m_cablesIn[11][16] ;
    output \m_cablesIn[12][16] ;
    output \m_cablesIn[12][17] ;
    input \B_int[13] ;
    input \m_cablesIn[11][13] ;
    input \B_int[14] ;
    input \m_cablesIn[11][14] ;
    output \m_cablesIn[12][14] ;
    output \m_cablesIn[12][15] ;
    input \B_int[11] ;
    input \m_cablesIn[11][11] ;
    input \B_int[12] ;
    input \m_cablesIn[11][12] ;
    output \m_cablesIn[12][12] ;
    output \m_cablesIn[12][13] ;
    input \B_int[9] ;
    input \m_cablesIn[11][9] ;
    input \B_int[10] ;
    input \m_cablesIn[11][10] ;
    output \m_cablesIn[12][10] ;
    output \m_cablesIn[12][11] ;
    input \B_int[7] ;
    input \m_cablesIn[11][7] ;
    input \B_int[8] ;
    input \m_cablesIn[11][8] ;
    output \m_cablesIn[12][8] ;
    output \m_cablesIn[12][9] ;
    input \B_int[5] ;
    input \m_cablesIn[11][5] ;
    input \B_int[6] ;
    input \m_cablesIn[11][6] ;
    output \m_cablesIn[12][6] ;
    output \m_cablesIn[12][7] ;
    input \B_int[3] ;
    input \m_cablesIn[11][3] ;
    input \B_int[4] ;
    input \m_cablesIn[11][4] ;
    output \m_cablesIn[12][4] ;
    output \m_cablesIn[12][5] ;
    input \B_int[1] ;
    input \m_cablesIn[11][1] ;
    input \B_int[2] ;
    input \m_cablesIn[11][2] ;
    output \m_cablesIn[12][2] ;
    output \m_cablesIn[12][3] ;
    input \B_int[0] ;
    input \frac_div[16] ;
    output \m_cablesIn[12][1] ;
    
    
    wire n62386, n62385, n62384, n62383, n62382, n62381, n62380, 
        n62379, n62378, n62377, n62376, n62375;
    
    CCU2D add_3381_25 (.A0(\m_cablesIn[11][23] ), .B0(\QQ_in[11][10] ), 
          .C0(GND_net), .D0(GND_net), .A1(\m_cablesIn[11][24] ), .B1(\QQ_in[11][10] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62386), .S0(\m_cablesIn[12][24] ), 
          .S1(\QQ_in[12][11] ));
    defparam add_3381_25.INIT0 = 16'h5666;
    defparam add_3381_25.INIT1 = 16'h5999;
    defparam add_3381_25.INJECT1_0 = "NO";
    defparam add_3381_25.INJECT1_1 = "NO";
    CCU2D add_3381_23 (.A0(\B_int[21] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][22] ), 
          .D1(GND_net), .CIN(n62385), .COUT(n62386), .S0(\m_cablesIn[12][22] ), 
          .S1(\m_cablesIn[12][23] ));
    defparam add_3381_23.INIT0 = 16'h6969;
    defparam add_3381_23.INIT1 = 16'h6969;
    defparam add_3381_23.INJECT1_0 = "NO";
    defparam add_3381_23.INJECT1_1 = "NO";
    CCU2D add_3381_21 (.A0(\B_int[19] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][20] ), 
          .D1(GND_net), .CIN(n62384), .COUT(n62385), .S0(\m_cablesIn[12][20] ), 
          .S1(\m_cablesIn[12][21] ));
    defparam add_3381_21.INIT0 = 16'h6969;
    defparam add_3381_21.INIT1 = 16'h6969;
    defparam add_3381_21.INJECT1_0 = "NO";
    defparam add_3381_21.INJECT1_1 = "NO";
    CCU2D add_3381_19 (.A0(\B_int[17] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][18] ), 
          .D1(GND_net), .CIN(n62383), .COUT(n62384), .S0(\m_cablesIn[12][18] ), 
          .S1(\m_cablesIn[12][19] ));
    defparam add_3381_19.INIT0 = 16'h6969;
    defparam add_3381_19.INIT1 = 16'h6969;
    defparam add_3381_19.INJECT1_0 = "NO";
    defparam add_3381_19.INJECT1_1 = "NO";
    CCU2D add_3381_17 (.A0(\B_int[15] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][16] ), 
          .D1(GND_net), .CIN(n62382), .COUT(n62383), .S0(\m_cablesIn[12][16] ), 
          .S1(\m_cablesIn[12][17] ));
    defparam add_3381_17.INIT0 = 16'h6969;
    defparam add_3381_17.INIT1 = 16'h6969;
    defparam add_3381_17.INJECT1_0 = "NO";
    defparam add_3381_17.INJECT1_1 = "NO";
    CCU2D add_3381_15 (.A0(\B_int[13] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][14] ), 
          .D1(GND_net), .CIN(n62381), .COUT(n62382), .S0(\m_cablesIn[12][14] ), 
          .S1(\m_cablesIn[12][15] ));
    defparam add_3381_15.INIT0 = 16'h6969;
    defparam add_3381_15.INIT1 = 16'h6969;
    defparam add_3381_15.INJECT1_0 = "NO";
    defparam add_3381_15.INJECT1_1 = "NO";
    CCU2D add_3381_13 (.A0(\B_int[11] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][12] ), 
          .D1(GND_net), .CIN(n62380), .COUT(n62381), .S0(\m_cablesIn[12][12] ), 
          .S1(\m_cablesIn[12][13] ));
    defparam add_3381_13.INIT0 = 16'h6969;
    defparam add_3381_13.INIT1 = 16'h6969;
    defparam add_3381_13.INJECT1_0 = "NO";
    defparam add_3381_13.INJECT1_1 = "NO";
    CCU2D add_3381_11 (.A0(\B_int[9] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][10] ), 
          .D1(GND_net), .CIN(n62379), .COUT(n62380), .S0(\m_cablesIn[12][10] ), 
          .S1(\m_cablesIn[12][11] ));
    defparam add_3381_11.INIT0 = 16'h6969;
    defparam add_3381_11.INIT1 = 16'h6969;
    defparam add_3381_11.INJECT1_0 = "NO";
    defparam add_3381_11.INJECT1_1 = "NO";
    CCU2D add_3381_9 (.A0(\B_int[7] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][8] ), 
          .D1(GND_net), .CIN(n62378), .COUT(n62379), .S0(\m_cablesIn[12][8] ), 
          .S1(\m_cablesIn[12][9] ));
    defparam add_3381_9.INIT0 = 16'h6969;
    defparam add_3381_9.INIT1 = 16'h6969;
    defparam add_3381_9.INJECT1_0 = "NO";
    defparam add_3381_9.INJECT1_1 = "NO";
    CCU2D add_3381_7 (.A0(\B_int[5] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][6] ), 
          .D1(GND_net), .CIN(n62377), .COUT(n62378), .S0(\m_cablesIn[12][6] ), 
          .S1(\m_cablesIn[12][7] ));
    defparam add_3381_7.INIT0 = 16'h6969;
    defparam add_3381_7.INIT1 = 16'h6969;
    defparam add_3381_7.INJECT1_0 = "NO";
    defparam add_3381_7.INJECT1_1 = "NO";
    CCU2D add_3381_5 (.A0(\B_int[3] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][4] ), 
          .D1(GND_net), .CIN(n62376), .COUT(n62377), .S0(\m_cablesIn[12][4] ), 
          .S1(\m_cablesIn[12][5] ));
    defparam add_3381_5.INIT0 = 16'h6969;
    defparam add_3381_5.INIT1 = 16'h6969;
    defparam add_3381_5.INJECT1_0 = "NO";
    defparam add_3381_5.INJECT1_1 = "NO";
    CCU2D add_3381_3 (.A0(\B_int[1] ), .B0(\QQ_in[11][10] ), .C0(\m_cablesIn[11][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[11][10] ), .C1(\m_cablesIn[11][2] ), 
          .D1(GND_net), .CIN(n62375), .COUT(n62376), .S0(\m_cablesIn[12][2] ), 
          .S1(\m_cablesIn[12][3] ));
    defparam add_3381_3.INIT0 = 16'h6969;
    defparam add_3381_3.INIT1 = 16'h6969;
    defparam add_3381_3.INJECT1_0 = "NO";
    defparam add_3381_3.INJECT1_1 = "NO";
    CCU2D add_3381_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[11][10] ), .C1(\frac_div[16] ), 
          .D1(GND_net), .COUT(n62375), .S1(\m_cablesIn[12][1] ));
    defparam add_3381_1.INIT0 = 16'hF000;
    defparam add_3381_1.INIT1 = 16'h6969;
    defparam add_3381_1.INJECT1_0 = "NO";
    defparam add_3381_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U23 
//

module \a_s(24)_U23  (\m_cablesIn[10][23] , \QQ_in[10][9] , GND_net, \m_cablesIn[10][24] , 
            \m_cablesIn[11][24] , \QQ_in[11][10] , \B_int[21] , \m_cablesIn[10][21] , 
            \B_int[22] , \m_cablesIn[10][22] , \m_cablesIn[11][22] , \m_cablesIn[11][23] , 
            \B_int[19] , \m_cablesIn[10][19] , \B_int[20] , \m_cablesIn[10][20] , 
            \m_cablesIn[11][20] , \m_cablesIn[11][21] , \B_int[17] , \m_cablesIn[10][17] , 
            \B_int[18] , \m_cablesIn[10][18] , \m_cablesIn[11][18] , \m_cablesIn[11][19] , 
            \B_int[15] , \m_cablesIn[10][15] , \B_int[16] , \m_cablesIn[10][16] , 
            \m_cablesIn[11][16] , \m_cablesIn[11][17] , \B_int[13] , \m_cablesIn[10][13] , 
            \B_int[14] , \m_cablesIn[10][14] , \m_cablesIn[11][14] , \m_cablesIn[11][15] , 
            \B_int[11] , \m_cablesIn[10][11] , \B_int[12] , \m_cablesIn[10][12] , 
            \m_cablesIn[11][12] , \m_cablesIn[11][13] , \B_int[9] , \m_cablesIn[10][9] , 
            \B_int[10] , \m_cablesIn[10][10] , \m_cablesIn[11][10] , \m_cablesIn[11][11] , 
            \B_int[7] , \m_cablesIn[10][7] , \B_int[8] , \m_cablesIn[10][8] , 
            \m_cablesIn[11][8] , \m_cablesIn[11][9] , \B_int[5] , \m_cablesIn[10][5] , 
            \B_int[6] , \m_cablesIn[10][6] , \m_cablesIn[11][6] , \m_cablesIn[11][7] , 
            \B_int[3] , \m_cablesIn[10][3] , \B_int[4] , \m_cablesIn[10][4] , 
            \m_cablesIn[11][4] , \m_cablesIn[11][5] , \B_int[1] , \m_cablesIn[10][1] , 
            \B_int[2] , \m_cablesIn[10][2] , \m_cablesIn[11][2] , \m_cablesIn[11][3] , 
            \B_int[0] , \frac_div[17] , \m_cablesIn[11][1] );
    input \m_cablesIn[10][23] ;
    input \QQ_in[10][9] ;
    input GND_net;
    input \m_cablesIn[10][24] ;
    output \m_cablesIn[11][24] ;
    output \QQ_in[11][10] ;
    input \B_int[21] ;
    input \m_cablesIn[10][21] ;
    input \B_int[22] ;
    input \m_cablesIn[10][22] ;
    output \m_cablesIn[11][22] ;
    output \m_cablesIn[11][23] ;
    input \B_int[19] ;
    input \m_cablesIn[10][19] ;
    input \B_int[20] ;
    input \m_cablesIn[10][20] ;
    output \m_cablesIn[11][20] ;
    output \m_cablesIn[11][21] ;
    input \B_int[17] ;
    input \m_cablesIn[10][17] ;
    input \B_int[18] ;
    input \m_cablesIn[10][18] ;
    output \m_cablesIn[11][18] ;
    output \m_cablesIn[11][19] ;
    input \B_int[15] ;
    input \m_cablesIn[10][15] ;
    input \B_int[16] ;
    input \m_cablesIn[10][16] ;
    output \m_cablesIn[11][16] ;
    output \m_cablesIn[11][17] ;
    input \B_int[13] ;
    input \m_cablesIn[10][13] ;
    input \B_int[14] ;
    input \m_cablesIn[10][14] ;
    output \m_cablesIn[11][14] ;
    output \m_cablesIn[11][15] ;
    input \B_int[11] ;
    input \m_cablesIn[10][11] ;
    input \B_int[12] ;
    input \m_cablesIn[10][12] ;
    output \m_cablesIn[11][12] ;
    output \m_cablesIn[11][13] ;
    input \B_int[9] ;
    input \m_cablesIn[10][9] ;
    input \B_int[10] ;
    input \m_cablesIn[10][10] ;
    output \m_cablesIn[11][10] ;
    output \m_cablesIn[11][11] ;
    input \B_int[7] ;
    input \m_cablesIn[10][7] ;
    input \B_int[8] ;
    input \m_cablesIn[10][8] ;
    output \m_cablesIn[11][8] ;
    output \m_cablesIn[11][9] ;
    input \B_int[5] ;
    input \m_cablesIn[10][5] ;
    input \B_int[6] ;
    input \m_cablesIn[10][6] ;
    output \m_cablesIn[11][6] ;
    output \m_cablesIn[11][7] ;
    input \B_int[3] ;
    input \m_cablesIn[10][3] ;
    input \B_int[4] ;
    input \m_cablesIn[10][4] ;
    output \m_cablesIn[11][4] ;
    output \m_cablesIn[11][5] ;
    input \B_int[1] ;
    input \m_cablesIn[10][1] ;
    input \B_int[2] ;
    input \m_cablesIn[10][2] ;
    output \m_cablesIn[11][2] ;
    output \m_cablesIn[11][3] ;
    input \B_int[0] ;
    input \frac_div[17] ;
    output \m_cablesIn[11][1] ;
    
    
    wire n62399, n62398, n62397, n62396, n62395, n62394, n62393, 
        n62392, n62391, n62390, n62389, n62388;
    
    CCU2D add_3355_25 (.A0(\m_cablesIn[10][23] ), .B0(\QQ_in[10][9] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[10][24] ), .B1(\QQ_in[10][9] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62399), .S0(\m_cablesIn[11][24] ), 
          .S1(\QQ_in[11][10] ));
    defparam add_3355_25.INIT0 = 16'h5666;
    defparam add_3355_25.INIT1 = 16'h5999;
    defparam add_3355_25.INJECT1_0 = "NO";
    defparam add_3355_25.INJECT1_1 = "NO";
    CCU2D add_3355_23 (.A0(\B_int[21] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][22] ), 
          .D1(GND_net), .CIN(n62398), .COUT(n62399), .S0(\m_cablesIn[11][22] ), 
          .S1(\m_cablesIn[11][23] ));
    defparam add_3355_23.INIT0 = 16'h6969;
    defparam add_3355_23.INIT1 = 16'h6969;
    defparam add_3355_23.INJECT1_0 = "NO";
    defparam add_3355_23.INJECT1_1 = "NO";
    CCU2D add_3355_21 (.A0(\B_int[19] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][20] ), 
          .D1(GND_net), .CIN(n62397), .COUT(n62398), .S0(\m_cablesIn[11][20] ), 
          .S1(\m_cablesIn[11][21] ));
    defparam add_3355_21.INIT0 = 16'h6969;
    defparam add_3355_21.INIT1 = 16'h6969;
    defparam add_3355_21.INJECT1_0 = "NO";
    defparam add_3355_21.INJECT1_1 = "NO";
    CCU2D add_3355_19 (.A0(\B_int[17] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][18] ), 
          .D1(GND_net), .CIN(n62396), .COUT(n62397), .S0(\m_cablesIn[11][18] ), 
          .S1(\m_cablesIn[11][19] ));
    defparam add_3355_19.INIT0 = 16'h6969;
    defparam add_3355_19.INIT1 = 16'h6969;
    defparam add_3355_19.INJECT1_0 = "NO";
    defparam add_3355_19.INJECT1_1 = "NO";
    CCU2D add_3355_17 (.A0(\B_int[15] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][16] ), 
          .D1(GND_net), .CIN(n62395), .COUT(n62396), .S0(\m_cablesIn[11][16] ), 
          .S1(\m_cablesIn[11][17] ));
    defparam add_3355_17.INIT0 = 16'h6969;
    defparam add_3355_17.INIT1 = 16'h6969;
    defparam add_3355_17.INJECT1_0 = "NO";
    defparam add_3355_17.INJECT1_1 = "NO";
    CCU2D add_3355_15 (.A0(\B_int[13] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][14] ), 
          .D1(GND_net), .CIN(n62394), .COUT(n62395), .S0(\m_cablesIn[11][14] ), 
          .S1(\m_cablesIn[11][15] ));
    defparam add_3355_15.INIT0 = 16'h6969;
    defparam add_3355_15.INIT1 = 16'h6969;
    defparam add_3355_15.INJECT1_0 = "NO";
    defparam add_3355_15.INJECT1_1 = "NO";
    CCU2D add_3355_13 (.A0(\B_int[11] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][12] ), 
          .D1(GND_net), .CIN(n62393), .COUT(n62394), .S0(\m_cablesIn[11][12] ), 
          .S1(\m_cablesIn[11][13] ));
    defparam add_3355_13.INIT0 = 16'h6969;
    defparam add_3355_13.INIT1 = 16'h6969;
    defparam add_3355_13.INJECT1_0 = "NO";
    defparam add_3355_13.INJECT1_1 = "NO";
    CCU2D add_3355_11 (.A0(\B_int[9] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][10] ), 
          .D1(GND_net), .CIN(n62392), .COUT(n62393), .S0(\m_cablesIn[11][10] ), 
          .S1(\m_cablesIn[11][11] ));
    defparam add_3355_11.INIT0 = 16'h6969;
    defparam add_3355_11.INIT1 = 16'h6969;
    defparam add_3355_11.INJECT1_0 = "NO";
    defparam add_3355_11.INJECT1_1 = "NO";
    CCU2D add_3355_9 (.A0(\B_int[7] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][8] ), 
          .D1(GND_net), .CIN(n62391), .COUT(n62392), .S0(\m_cablesIn[11][8] ), 
          .S1(\m_cablesIn[11][9] ));
    defparam add_3355_9.INIT0 = 16'h6969;
    defparam add_3355_9.INIT1 = 16'h6969;
    defparam add_3355_9.INJECT1_0 = "NO";
    defparam add_3355_9.INJECT1_1 = "NO";
    CCU2D add_3355_7 (.A0(\B_int[5] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][6] ), 
          .D1(GND_net), .CIN(n62390), .COUT(n62391), .S0(\m_cablesIn[11][6] ), 
          .S1(\m_cablesIn[11][7] ));
    defparam add_3355_7.INIT0 = 16'h6969;
    defparam add_3355_7.INIT1 = 16'h6969;
    defparam add_3355_7.INJECT1_0 = "NO";
    defparam add_3355_7.INJECT1_1 = "NO";
    CCU2D add_3355_5 (.A0(\B_int[3] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][4] ), 
          .D1(GND_net), .CIN(n62389), .COUT(n62390), .S0(\m_cablesIn[11][4] ), 
          .S1(\m_cablesIn[11][5] ));
    defparam add_3355_5.INIT0 = 16'h6969;
    defparam add_3355_5.INIT1 = 16'h6969;
    defparam add_3355_5.INJECT1_0 = "NO";
    defparam add_3355_5.INJECT1_1 = "NO";
    CCU2D add_3355_3 (.A0(\B_int[1] ), .B0(\QQ_in[10][9] ), .C0(\m_cablesIn[10][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[10][9] ), .C1(\m_cablesIn[10][2] ), 
          .D1(GND_net), .CIN(n62388), .COUT(n62389), .S0(\m_cablesIn[11][2] ), 
          .S1(\m_cablesIn[11][3] ));
    defparam add_3355_3.INIT0 = 16'h6969;
    defparam add_3355_3.INIT1 = 16'h6969;
    defparam add_3355_3.INJECT1_0 = "NO";
    defparam add_3355_3.INJECT1_1 = "NO";
    CCU2D add_3355_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[10][9] ), .C1(\frac_div[17] ), .D1(GND_net), 
          .COUT(n62388), .S1(\m_cablesIn[11][1] ));
    defparam add_3355_1.INIT0 = 16'hF000;
    defparam add_3355_1.INIT1 = 16'h6969;
    defparam add_3355_1.INJECT1_0 = "NO";
    defparam add_3355_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \a_s(24)_U24 
//

module \a_s(24)_U24  (\m_cablesIn[9][23] , \QQ_in[9][8] , GND_net, \m_cablesIn[9][24] , 
            \m_cablesIn[10][24] , \QQ_in[10][9] , \B_int[21] , \m_cablesIn[9][21] , 
            \B_int[22] , \m_cablesIn[9][22] , \m_cablesIn[10][22] , \m_cablesIn[10][23] , 
            \B_int[19] , \m_cablesIn[9][19] , \B_int[20] , \m_cablesIn[9][20] , 
            \m_cablesIn[10][20] , \m_cablesIn[10][21] , \B_int[17] , \m_cablesIn[9][17] , 
            \B_int[18] , \m_cablesIn[9][18] , \m_cablesIn[10][18] , \m_cablesIn[10][19] , 
            \B_int[15] , \m_cablesIn[9][15] , \B_int[16] , \m_cablesIn[9][16] , 
            \m_cablesIn[10][16] , \m_cablesIn[10][17] , \B_int[13] , \m_cablesIn[9][13] , 
            \B_int[14] , \m_cablesIn[9][14] , \m_cablesIn[10][14] , \m_cablesIn[10][15] , 
            \B_int[11] , \m_cablesIn[9][11] , \B_int[12] , \m_cablesIn[9][12] , 
            \m_cablesIn[10][12] , \m_cablesIn[10][13] , \B_int[9] , \m_cablesIn[9][9] , 
            \B_int[10] , \m_cablesIn[9][10] , \m_cablesIn[10][10] , \m_cablesIn[10][11] , 
            \B_int[7] , \m_cablesIn[9][7] , \B_int[8] , \m_cablesIn[9][8] , 
            \m_cablesIn[10][8] , \m_cablesIn[10][9] , \B_int[5] , \m_cablesIn[9][5] , 
            \B_int[6] , \m_cablesIn[9][6] , \m_cablesIn[10][6] , \m_cablesIn[10][7] , 
            \B_int[3] , \m_cablesIn[9][3] , \B_int[4] , \m_cablesIn[9][4] , 
            \m_cablesIn[10][4] , \m_cablesIn[10][5] , \B_int[1] , \m_cablesIn[9][1] , 
            \B_int[2] , \m_cablesIn[9][2] , \m_cablesIn[10][2] , \m_cablesIn[10][3] , 
            \B_int[0] , \frac_div[18] , \m_cablesIn[10][1] );
    input \m_cablesIn[9][23] ;
    input \QQ_in[9][8] ;
    input GND_net;
    input \m_cablesIn[9][24] ;
    output \m_cablesIn[10][24] ;
    output \QQ_in[10][9] ;
    input \B_int[21] ;
    input \m_cablesIn[9][21] ;
    input \B_int[22] ;
    input \m_cablesIn[9][22] ;
    output \m_cablesIn[10][22] ;
    output \m_cablesIn[10][23] ;
    input \B_int[19] ;
    input \m_cablesIn[9][19] ;
    input \B_int[20] ;
    input \m_cablesIn[9][20] ;
    output \m_cablesIn[10][20] ;
    output \m_cablesIn[10][21] ;
    input \B_int[17] ;
    input \m_cablesIn[9][17] ;
    input \B_int[18] ;
    input \m_cablesIn[9][18] ;
    output \m_cablesIn[10][18] ;
    output \m_cablesIn[10][19] ;
    input \B_int[15] ;
    input \m_cablesIn[9][15] ;
    input \B_int[16] ;
    input \m_cablesIn[9][16] ;
    output \m_cablesIn[10][16] ;
    output \m_cablesIn[10][17] ;
    input \B_int[13] ;
    input \m_cablesIn[9][13] ;
    input \B_int[14] ;
    input \m_cablesIn[9][14] ;
    output \m_cablesIn[10][14] ;
    output \m_cablesIn[10][15] ;
    input \B_int[11] ;
    input \m_cablesIn[9][11] ;
    input \B_int[12] ;
    input \m_cablesIn[9][12] ;
    output \m_cablesIn[10][12] ;
    output \m_cablesIn[10][13] ;
    input \B_int[9] ;
    input \m_cablesIn[9][9] ;
    input \B_int[10] ;
    input \m_cablesIn[9][10] ;
    output \m_cablesIn[10][10] ;
    output \m_cablesIn[10][11] ;
    input \B_int[7] ;
    input \m_cablesIn[9][7] ;
    input \B_int[8] ;
    input \m_cablesIn[9][8] ;
    output \m_cablesIn[10][8] ;
    output \m_cablesIn[10][9] ;
    input \B_int[5] ;
    input \m_cablesIn[9][5] ;
    input \B_int[6] ;
    input \m_cablesIn[9][6] ;
    output \m_cablesIn[10][6] ;
    output \m_cablesIn[10][7] ;
    input \B_int[3] ;
    input \m_cablesIn[9][3] ;
    input \B_int[4] ;
    input \m_cablesIn[9][4] ;
    output \m_cablesIn[10][4] ;
    output \m_cablesIn[10][5] ;
    input \B_int[1] ;
    input \m_cablesIn[9][1] ;
    input \B_int[2] ;
    input \m_cablesIn[9][2] ;
    output \m_cablesIn[10][2] ;
    output \m_cablesIn[10][3] ;
    input \B_int[0] ;
    input \frac_div[18] ;
    output \m_cablesIn[10][1] ;
    
    
    wire n62412, n62411, n62410, n62409, n62408, n62407, n62406, 
        n62405, n62404, n62403, n62402, n62401;
    
    CCU2D add_3329_25 (.A0(\m_cablesIn[9][23] ), .B0(\QQ_in[9][8] ), .C0(GND_net), 
          .D0(GND_net), .A1(\m_cablesIn[9][24] ), .B1(\QQ_in[9][8] ), 
          .C1(GND_net), .D1(GND_net), .CIN(n62412), .S0(\m_cablesIn[10][24] ), 
          .S1(\QQ_in[10][9] ));
    defparam add_3329_25.INIT0 = 16'h5666;
    defparam add_3329_25.INIT1 = 16'h5999;
    defparam add_3329_25.INJECT1_0 = "NO";
    defparam add_3329_25.INJECT1_1 = "NO";
    CCU2D add_3329_23 (.A0(\B_int[21] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][21] ), 
          .D0(GND_net), .A1(\B_int[22] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][22] ), 
          .D1(GND_net), .CIN(n62411), .COUT(n62412), .S0(\m_cablesIn[10][22] ), 
          .S1(\m_cablesIn[10][23] ));
    defparam add_3329_23.INIT0 = 16'h6969;
    defparam add_3329_23.INIT1 = 16'h6969;
    defparam add_3329_23.INJECT1_0 = "NO";
    defparam add_3329_23.INJECT1_1 = "NO";
    CCU2D add_3329_21 (.A0(\B_int[19] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][19] ), 
          .D0(GND_net), .A1(\B_int[20] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][20] ), 
          .D1(GND_net), .CIN(n62410), .COUT(n62411), .S0(\m_cablesIn[10][20] ), 
          .S1(\m_cablesIn[10][21] ));
    defparam add_3329_21.INIT0 = 16'h6969;
    defparam add_3329_21.INIT1 = 16'h6969;
    defparam add_3329_21.INJECT1_0 = "NO";
    defparam add_3329_21.INJECT1_1 = "NO";
    CCU2D add_3329_19 (.A0(\B_int[17] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][17] ), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][18] ), 
          .D1(GND_net), .CIN(n62409), .COUT(n62410), .S0(\m_cablesIn[10][18] ), 
          .S1(\m_cablesIn[10][19] ));
    defparam add_3329_19.INIT0 = 16'h6969;
    defparam add_3329_19.INIT1 = 16'h6969;
    defparam add_3329_19.INJECT1_0 = "NO";
    defparam add_3329_19.INJECT1_1 = "NO";
    CCU2D add_3329_17 (.A0(\B_int[15] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][15] ), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][16] ), 
          .D1(GND_net), .CIN(n62408), .COUT(n62409), .S0(\m_cablesIn[10][16] ), 
          .S1(\m_cablesIn[10][17] ));
    defparam add_3329_17.INIT0 = 16'h6969;
    defparam add_3329_17.INIT1 = 16'h6969;
    defparam add_3329_17.INJECT1_0 = "NO";
    defparam add_3329_17.INJECT1_1 = "NO";
    CCU2D add_3329_15 (.A0(\B_int[13] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][13] ), 
          .D0(GND_net), .A1(\B_int[14] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][14] ), 
          .D1(GND_net), .CIN(n62407), .COUT(n62408), .S0(\m_cablesIn[10][14] ), 
          .S1(\m_cablesIn[10][15] ));
    defparam add_3329_15.INIT0 = 16'h6969;
    defparam add_3329_15.INIT1 = 16'h6969;
    defparam add_3329_15.INJECT1_0 = "NO";
    defparam add_3329_15.INJECT1_1 = "NO";
    CCU2D add_3329_13 (.A0(\B_int[11] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][11] ), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][12] ), 
          .D1(GND_net), .CIN(n62406), .COUT(n62407), .S0(\m_cablesIn[10][12] ), 
          .S1(\m_cablesIn[10][13] ));
    defparam add_3329_13.INIT0 = 16'h6969;
    defparam add_3329_13.INIT1 = 16'h6969;
    defparam add_3329_13.INJECT1_0 = "NO";
    defparam add_3329_13.INJECT1_1 = "NO";
    CCU2D add_3329_11 (.A0(\B_int[9] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][9] ), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][10] ), 
          .D1(GND_net), .CIN(n62405), .COUT(n62406), .S0(\m_cablesIn[10][10] ), 
          .S1(\m_cablesIn[10][11] ));
    defparam add_3329_11.INIT0 = 16'h6969;
    defparam add_3329_11.INIT1 = 16'h6969;
    defparam add_3329_11.INJECT1_0 = "NO";
    defparam add_3329_11.INJECT1_1 = "NO";
    CCU2D add_3329_9 (.A0(\B_int[7] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][7] ), 
          .D0(GND_net), .A1(\B_int[8] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][8] ), 
          .D1(GND_net), .CIN(n62404), .COUT(n62405), .S0(\m_cablesIn[10][8] ), 
          .S1(\m_cablesIn[10][9] ));
    defparam add_3329_9.INIT0 = 16'h6969;
    defparam add_3329_9.INIT1 = 16'h6969;
    defparam add_3329_9.INJECT1_0 = "NO";
    defparam add_3329_9.INJECT1_1 = "NO";
    CCU2D add_3329_7 (.A0(\B_int[5] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][5] ), 
          .D0(GND_net), .A1(\B_int[6] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][6] ), 
          .D1(GND_net), .CIN(n62403), .COUT(n62404), .S0(\m_cablesIn[10][6] ), 
          .S1(\m_cablesIn[10][7] ));
    defparam add_3329_7.INIT0 = 16'h6969;
    defparam add_3329_7.INIT1 = 16'h6969;
    defparam add_3329_7.INJECT1_0 = "NO";
    defparam add_3329_7.INJECT1_1 = "NO";
    CCU2D add_3329_5 (.A0(\B_int[3] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][3] ), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][4] ), 
          .D1(GND_net), .CIN(n62402), .COUT(n62403), .S0(\m_cablesIn[10][4] ), 
          .S1(\m_cablesIn[10][5] ));
    defparam add_3329_5.INIT0 = 16'h6969;
    defparam add_3329_5.INIT1 = 16'h6969;
    defparam add_3329_5.INJECT1_0 = "NO";
    defparam add_3329_5.INJECT1_1 = "NO";
    CCU2D add_3329_3 (.A0(\B_int[1] ), .B0(\QQ_in[9][8] ), .C0(\m_cablesIn[9][1] ), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\QQ_in[9][8] ), .C1(\m_cablesIn[9][2] ), 
          .D1(GND_net), .CIN(n62401), .COUT(n62402), .S0(\m_cablesIn[10][2] ), 
          .S1(\m_cablesIn[10][3] ));
    defparam add_3329_3.INIT0 = 16'h6969;
    defparam add_3329_3.INIT1 = 16'h6969;
    defparam add_3329_3.INJECT1_0 = "NO";
    defparam add_3329_3.INJECT1_1 = "NO";
    CCU2D add_3329_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\B_int[0] ), .B1(\QQ_in[9][8] ), .C1(\frac_div[18] ), .D1(GND_net), 
          .COUT(n62401), .S1(\m_cablesIn[10][1] ));
    defparam add_3329_1.INIT0 = 16'hF000;
    defparam add_3329_1.INIT1 = 16'h6969;
    defparam add_3329_1.INJECT1_0 = "NO";
    defparam add_3329_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \fp_add(32,24,8)_U28 
//

module \fp_add(32,24,8)_U28  (add_c, clock, n73804, \A_int[11] , \B_int[11] , 
            \A_int[10] , \B_int[10] , \A_int[13] , \B_int[13] , \A_int[12] , 
            \B_int[12] , add_ce, \A_int[17] , \B_int[17] , alu_b, 
            \A_int[16] , \B_int[16] , alu_a, \A_int[18] , \B_int[18] , 
            GND_net, \A_int[2] , \B_int[2] , \B_int[3] , \A_int[9] , 
            \A_int[7] , \A_int[4] , \A_int[3] , \B_int[9] , \B_int[7] , 
            \B_int[4] , diffExpAB, add_enable, \diffExp[4] , n73803, 
            n70835, n70834, n70833, \efectFracB[21] , \efectFracB[20] , 
            \efectFracB[19] , \efectFracB[15] , \efectFracB[16] , n19214, 
            n28, n70771, n9, \efectFracB[14] , \efectFracB[7] , \efectFracB[5] , 
            \efectFracB[12] , n70820, \efectFracB[13] , n27, n70740, 
            n55);
    output [31:0]add_c;
    input clock;
    input n73804;
    output \A_int[11] ;
    output \B_int[11] ;
    output \A_int[10] ;
    output \B_int[10] ;
    output \A_int[13] ;
    output \B_int[13] ;
    output \A_int[12] ;
    output \B_int[12] ;
    input add_ce;
    output \A_int[17] ;
    output \B_int[17] ;
    input [31:0]alu_b;
    output \A_int[16] ;
    output \B_int[16] ;
    input [31:0]alu_a;
    output \A_int[18] ;
    output \B_int[18] ;
    input GND_net;
    output \A_int[2] ;
    output \B_int[2] ;
    output \B_int[3] ;
    output \A_int[9] ;
    output \A_int[7] ;
    output \A_int[4] ;
    output \A_int[3] ;
    output \B_int[9] ;
    output \B_int[7] ;
    output \B_int[4] ;
    output [8:0]diffExpAB;
    input add_enable;
    output \diffExp[4] ;
    input n73803;
    output n70835;
    output n70834;
    output n70833;
    input \efectFracB[21] ;
    input \efectFracB[20] ;
    input \efectFracB[19] ;
    input \efectFracB[15] ;
    input \efectFracB[16] ;
    input n19214;
    input n28;
    input n70771;
    input n9;
    input \efectFracB[14] ;
    input \efectFracB[7] ;
    input \efectFracB[5] ;
    input \efectFracB[12] ;
    input n70820;
    input \efectFracB[13] ;
    input n27;
    input n70740;
    input n55;
    
    wire [27:0]addSubAB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(69[18:26])
    wire [27:0]subBAExpEq;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(73[11:21])
    wire [31:0]A_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(54[11:16])
    wire [31:0]B_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(55[11:16])
    wire [31:0]FP_Z_int;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(106[11:19])
    wire [22:0]frac_Norm2;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(98[11:21])
    wire [27:0]frac;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(97[11:15])
    wire [27:0]frac_add_Norm1;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(70[11:25])
    wire [4:0]leadZerosBin;   // c:/users/yisong/documents/new/mlp/fp_leading_zeros_and_shift.vhd(25[11:23])
    wire [27:0]fracAlign_int;   // c:/users/yisong/documents/new/mlp/right_shifter.vhd(21[11:24])
    wire [8:0]efectExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(65[11:19])
    wire expB_FF;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(56[20:27])
    wire [8:0]diffExpBA;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[22:31])
    wire sign;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(75[11:15])
    wire isSUB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(71[11:16])
    wire [27:0]frac_sub_Norm1;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(74[11:25])
    wire [27:0]frac_Norm1;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(97[17:27])
    wire [8:0]diffExpAB_c;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[11:20])
    wire expA_FF;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(56[11:18])
    wire [27:0]efectFracB_align;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(67[35:51])
    wire [8:0]diffExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[33:40])
    
    wire n70733;
    wire [27:0]n451;
    
    wire n24122;
    wire [22:0]n10673;
    
    wire n70737;
    wire [27:0]n480;
    
    wire n770, n769, n768, n767, n766, n70739, n70613, n765, 
        n764, n763, n10, n70707, n70706, n17;
    wire [27:0]n330;
    
    wire n18, n70714, n15, n70865, n448, n7, n21713, n21711, 
        n21685, n21687, n21675, n21661, n21663, n21659, n21677, 
        n21657, n21671, n21667, n21653, n21655, n21665, n21641, 
        n21647, n21681, n62965, n53, n23602;
    wire [7:0]n8360;
    
    wire n70784, n40687, n66234, n731, n14, n66206, n9_c, n14_adj_418, 
        n10_adj_419, n67677, n61859, n60992, n28_c, n61858, n70715, 
        n31, n24, n70805, n36, n29, n26, n70703, n34, n66182, 
        n38, n25, n41758, n61857, n61856, n70726, n38_adj_420, 
        n24_adj_421, n36_adj_422, n42, n32, n31_adj_423, n70641, 
        n39, n70643, n70638;
    wire [27:0]n243;
    
    wire n40, n19140;
    wire [27:0]n272;
    
    wire n60991, n4, n44, n70636, n70637, n40002, n31_adj_424, 
        n66192, n28_adj_425, n38_adj_426, n24_adj_427, n10_adj_428, 
        n36_adj_429, n42_adj_430, n19142, n32_adj_431, n40_adj_432, 
        n44_adj_433, n31_adj_434, n19138, n66653, n70633, n14_adj_435, 
        n73795, n21808, n66558, n19, n63661, n63665, n61531, n61530, 
        n61529, n61528, n61527, n61526, n61525, n61524, n61523, 
        n61522, n61521, n61520, n17318, n61518, n62218, n62217, 
        n21643, n66178, n62216, n21651, n21645, n14_adj_436, n13, 
        n62215, n62214, n21679, n62213, n61517, n62212, n62211, 
        n61516, n62210, n21669, n61515, n62209, n62208, n62207, 
        n62206, n62205, n61513, n37, n39_adj_437, n34_adj_438, n61512, 
        n41, n30, n45, n4_adj_439, n44_adj_440, n33, n48, n43, 
        n574, n61511, n61510, n61509, n61508, n61507, n61506, 
        n61505, n61504, n61503, n13_adj_441, n41510, n41506, n41508, 
        n41778, n16, n15_adj_442, n70777, n41588, n15_adj_443, n70743, 
        n66914, n66904, n70832, n22565, n61613, n61612, n61611, 
        n70623, n61610;
    
    LUT4 mux_51_i13_3_lut (.A(addSubAB[12]), .B(subBAExpEq[12]), .C(n70733), 
         .Z(n451[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i13_3_lut.init = 16'hcaca;
    FD1P3IX FP_Z_i0_i19 (.D(n10673[19]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[19]));
    defparam FP_Z_i0_i19.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i20 (.D(n10673[20]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[20]));
    defparam FP_Z_i0_i20.GSR = "DISABLED";
    LUT4 mux_52_i12_3_lut (.A(A_int[8]), .B(B_int[8]), .C(n70737), .Z(n480[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i12_3_lut.init = 16'hacac;
    LUT4 mux_51_i12_3_lut (.A(addSubAB[11]), .B(subBAExpEq[11]), .C(n70733), 
         .Z(n451[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i12_3_lut.init = 16'hcaca;
    FD1P3IX FP_Z_i0_i21 (.D(n10673[21]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[21]));
    defparam FP_Z_i0_i21.GSR = "DISABLED";
    LUT4 mux_52_i15_3_lut (.A(\A_int[11] ), .B(\B_int[11] ), .C(n70737), 
         .Z(n480[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i15_3_lut.init = 16'hacac;
    LUT4 mux_51_i15_3_lut (.A(addSubAB[14]), .B(subBAExpEq[14]), .C(n70733), 
         .Z(n451[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i15_3_lut.init = 16'hcaca;
    FD1P3IX FP_Z_i0_i22 (.D(n10673[22]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[22]));
    defparam FP_Z_i0_i22.GSR = "DISABLED";
    LUT4 mux_52_i14_3_lut (.A(\A_int[10] ), .B(\B_int[10] ), .C(n70737), 
         .Z(n480[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i14_3_lut.init = 16'hacac;
    LUT4 mux_51_i14_3_lut (.A(addSubAB[13]), .B(subBAExpEq[13]), .C(n70733), 
         .Z(n451[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i14_3_lut.init = 16'hcaca;
    LUT4 mux_52_i17_3_lut (.A(\A_int[13] ), .B(\B_int[13] ), .C(n70737), 
         .Z(n480[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i17_3_lut.init = 16'hacac;
    FD1P3JX FP_Z_i0_i23 (.D(n770), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[23]));
    defparam FP_Z_i0_i23.GSR = "DISABLED";
    LUT4 mux_51_i17_3_lut (.A(addSubAB[16]), .B(subBAExpEq[16]), .C(n70733), 
         .Z(n451[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i17_3_lut.init = 16'hcaca;
    LUT4 mux_52_i16_3_lut (.A(\A_int[12] ), .B(\B_int[12] ), .C(n70737), 
         .Z(n480[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i16_3_lut.init = 16'hacac;
    LUT4 mux_51_i16_3_lut (.A(addSubAB[15]), .B(subBAExpEq[15]), .C(n70733), 
         .Z(n451[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i16_3_lut.init = 16'hcaca;
    LUT4 mux_52_i19_3_lut (.A(A_int[15]), .B(B_int[15]), .C(n70737), .Z(n480[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i19_3_lut.init = 16'hacac;
    FD1P3JX FP_Z_i0_i24 (.D(n769), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[24]));
    defparam FP_Z_i0_i24.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i15 (.D(n10673[15]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[15]));
    defparam FP_Z_i0_i15.GSR = "DISABLED";
    LUT4 mux_51_i19_3_lut (.A(addSubAB[18]), .B(subBAExpEq[18]), .C(n70733), 
         .Z(n451[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i19_3_lut.init = 16'hcaca;
    LUT4 mux_52_i18_3_lut (.A(A_int[14]), .B(B_int[14]), .C(n70737), .Z(n480[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i18_3_lut.init = 16'hacac;
    FD1P3JX FP_Z_i0_i25 (.D(n768), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[25]));
    defparam FP_Z_i0_i25.GSR = "DISABLED";
    LUT4 mux_51_i18_3_lut (.A(addSubAB[17]), .B(subBAExpEq[17]), .C(n70733), 
         .Z(n451[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i18_3_lut.init = 16'hcaca;
    LUT4 mux_52_i21_3_lut (.A(\A_int[17] ), .B(\B_int[17] ), .C(n70737), 
         .Z(n480[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i21_3_lut.init = 16'hacac;
    LUT4 mux_51_i21_3_lut (.A(addSubAB[20]), .B(subBAExpEq[20]), .C(n70733), 
         .Z(n451[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i21_3_lut.init = 16'hcaca;
    FD1P3AX B_int_i0_i0 (.D(alu_b[0]), .SP(n73804), .CK(clock), .Q(B_int[0]));
    defparam B_int_i0_i0.GSR = "DISABLED";
    LUT4 mux_52_i20_3_lut (.A(\A_int[16] ), .B(\B_int[16] ), .C(n70737), 
         .Z(n480[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i20_3_lut.init = 16'hacac;
    FD1P3AX FP_Z_i0_i0 (.D(FP_Z_int[0]), .SP(n73804), .CK(clock), .Q(add_c[0]));
    defparam FP_Z_i0_i0.GSR = "DISABLED";
    FD1P3AX A_int_i0_i0 (.D(alu_a[0]), .SP(n73804), .CK(clock), .Q(A_int[0]));
    defparam A_int_i0_i0.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i16 (.D(n10673[16]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[16]));
    defparam FP_Z_i0_i16.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i26 (.D(n767), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[26]));
    defparam FP_Z_i0_i26.GSR = "DISABLED";
    LUT4 mux_51_i20_3_lut (.A(addSubAB[19]), .B(subBAExpEq[19]), .C(n70733), 
         .Z(n451[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i20_3_lut.init = 16'hcaca;
    LUT4 mux_52_i23_3_lut (.A(A_int[19]), .B(B_int[19]), .C(n70737), .Z(n480[22])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i23_3_lut.init = 16'hacac;
    FD1P3IX FP_Z_i0_i17 (.D(n10673[17]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[17]));
    defparam FP_Z_i0_i17.GSR = "DISABLED";
    LUT4 mux_51_i23_3_lut (.A(addSubAB[22]), .B(subBAExpEq[22]), .C(n70733), 
         .Z(n451[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i23_3_lut.init = 16'hcaca;
    LUT4 mux_52_i22_3_lut (.A(\A_int[18] ), .B(\B_int[18] ), .C(n70737), 
         .Z(n480[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i22_3_lut.init = 16'hacac;
    LUT4 mux_51_i22_3_lut (.A(addSubAB[21]), .B(subBAExpEq[21]), .C(n70733), 
         .Z(n451[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i22_3_lut.init = 16'hcaca;
    LUT4 mux_52_i25_3_lut (.A(A_int[21]), .B(B_int[21]), .C(n70737), .Z(n480[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i25_3_lut.init = 16'hacac;
    FD1P3JX FP_Z_i0_i27 (.D(n766), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[27]));
    defparam FP_Z_i0_i27.GSR = "DISABLED";
    LUT4 mux_51_i25_3_lut (.A(addSubAB[24]), .B(subBAExpEq[24]), .C(n70733), 
         .Z(n451[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i25_3_lut.init = 16'hcaca;
    FD1P3IX FP_Z_i0_i18 (.D(n10673[18]), .SP(n73804), .CD(n24122), .CK(clock), 
            .Q(add_c[18]));
    defparam FP_Z_i0_i18.GSR = "DISABLED";
    LUT4 mux_52_i24_3_lut (.A(A_int[20]), .B(B_int[20]), .C(n70737), .Z(n480[23])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i24_3_lut.init = 16'hacac;
    LUT4 mux_3773_i22_4_lut (.A(frac_Norm2[21]), .B(frac[24]), .C(n70739), 
         .D(n70613), .Z(n10673[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i22_4_lut.init = 16'hcac0;
    FD1P3JX FP_Z_i0_i28 (.D(n765), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[28]));
    defparam FP_Z_i0_i28.GSR = "DISABLED";
    LUT4 mux_51_i24_3_lut (.A(addSubAB[23]), .B(subBAExpEq[23]), .C(n70733), 
         .Z(n451[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i24_3_lut.init = 16'hcaca;
    LUT4 mux_52_i26_3_lut (.A(A_int[22]), .B(B_int[22]), .C(n70737), .Z(n480[25])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i26_3_lut.init = 16'hacac;
    LUT4 mux_51_i26_3_lut (.A(addSubAB[25]), .B(subBAExpEq[25]), .C(n70733), 
         .Z(n451[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i26_3_lut.init = 16'hcaca;
    FD1P3JX FP_Z_i0_i29 (.D(n764), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[29]));
    defparam FP_Z_i0_i29.GSR = "DISABLED";
    FD1P3JX FP_Z_i0_i30 (.D(n763), .SP(n73804), .PD(n24122), .CK(clock), 
            .Q(add_c[30]));
    defparam FP_Z_i0_i30.GSR = "DISABLED";
    LUT4 i2_2_lut (.A(B_int[25]), .B(B_int[27]), .Z(n10)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 mux_216_i4_3_lut (.A(n70707), .B(n70706), .C(frac[27]), .Z(frac_add_Norm1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i4_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(n17), .B(n330[2]), .C(leadZerosBin[2]), .Z(n18)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut.init = 16'h0808;
    LUT4 i1_4_lut (.A(n70707), .B(n70714), .C(n70706), .D(frac[27]), 
         .Z(n15)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i1_3_lut_rep_763_4_lut (.A(A_int[31]), .B(n70865), .C(n448), 
         .D(subBAExpEq[27]), .Z(n70733)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B+((D)+!C)))) */ ;
    defparam i1_3_lut_rep_763_4_lut.init = 16'h0090;
    LUT4 i1_3_lut_4_lut (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[4]), 
         .Z(n21713)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_764 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[3]), 
         .Z(n21711)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_764.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_765 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[6]), 
         .Z(n21685)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_765.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_766 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[5]), 
         .Z(n21687)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_766.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_767 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[8]), 
         .Z(n21675)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_767.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_768 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[7]), 
         .Z(n21661)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_768.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_769 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[10]), 
         .Z(n21663)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_769.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_770 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[9]), 
         .Z(n21659)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_770.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_771 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[12]), 
         .Z(n21677)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_771.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_772 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[14]), 
         .Z(n21657)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_772.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_773 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[13]), 
         .Z(n21671)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_773.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_774 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[16]), 
         .Z(n21667)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_774.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_775 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[15]), 
         .Z(n21653)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_775.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_776 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[18]), 
         .Z(n21655)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_776.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_777 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[17]), 
         .Z(n21665)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_777.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_778 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[22]), 
         .Z(n21641)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_778.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_779 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[20]), 
         .Z(n21647)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_779.init = 16'h6966;
    LUT4 i1_3_lut_4_lut_adj_780 (.A(A_int[31]), .B(n70865), .C(n7), .D(fracAlign_int[21]), 
         .Z(n21681)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_780.init = 16'h6966;
    LUT4 i28155_3_lut_rep_643_4_lut (.A(A_int[31]), .B(n70865), .C(n62965), 
         .D(n53), .Z(n70613)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B+(C (D)))) */ ;
    defparam i28155_3_lut_rep_643_4_lut.init = 16'hf666;
    LUT4 i11916_3_lut (.A(addSubAB[1]), .B(addSubAB[2]), .C(frac[27]), 
         .Z(n23602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11916_3_lut.init = 16'hcaca;
    LUT4 i114_4_lut (.A(n8360[3]), .B(n70784), .C(n70739), .D(n40687), 
         .Z(n767)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i114_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i17_4_lut (.A(frac_Norm2[16]), .B(frac[19]), .C(n70739), 
         .D(n70613), .Z(n10673[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i17_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i15_4_lut (.A(frac_Norm2[14]), .B(frac[17]), .C(n70739), 
         .D(n70613), .Z(n10673[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i15_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i14_4_lut (.A(frac_Norm2[13]), .B(frac[16]), .C(n70739), 
         .D(n70613), .Z(n10673[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i14_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i13_4_lut (.A(frac_Norm2[12]), .B(frac[15]), .C(n70739), 
         .D(n70613), .Z(n10673[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i13_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i12_4_lut (.A(frac_Norm2[11]), .B(frac[14]), .C(n70739), 
         .D(n70613), .Z(n10673[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i12_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i11_4_lut (.A(frac_Norm2[10]), .B(frac[13]), .C(n70739), 
         .D(n70613), .Z(n10673[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i11_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i10_4_lut (.A(frac_Norm2[9]), .B(frac[12]), .C(n70739), 
         .D(n70613), .Z(n10673[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i10_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i9_4_lut (.A(frac_Norm2[8]), .B(frac[11]), .C(n70739), 
         .D(n70613), .Z(n10673[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i9_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i8_4_lut (.A(frac_Norm2[7]), .B(frac[10]), .C(n70739), 
         .D(n70613), .Z(n10673[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i8_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i7_4_lut (.A(frac_Norm2[6]), .B(frac[9]), .C(n70739), 
         .D(n70613), .Z(n10673[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i7_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i6_4_lut (.A(frac_Norm2[5]), .B(frac[8]), .C(n70739), 
         .D(n70613), .Z(n10673[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i6_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i1_4_lut (.A(frac_Norm2[0]), .B(n70707), .C(n70739), 
         .D(n70613), .Z(n10673[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i1_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i5_4_lut (.A(frac_Norm2[4]), .B(frac[7]), .C(n70739), 
         .D(n70613), .Z(n10673[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i5_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut (.A(n10673[0]), .B(n66234), .C(n731), .Z(FP_Z_int[0])) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i1_3_lut.init = 16'hcece;
    LUT4 i6_4_lut (.A(B_int[26]), .B(B_int[24]), .C(B_int[28]), .D(B_int[30]), 
         .Z(n14)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i115_4_lut (.A(n8360[2]), .B(efectExp[2]), .C(n70739), .D(n40687), 
         .Z(n768)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i115_4_lut.init = 16'hcac0;
    LUT4 i7_4_lut (.A(B_int[23]), .B(n14), .C(n10), .D(B_int[29]), .Z(expB_FF)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'h8000;
    LUT4 mux_3773_i16_4_lut (.A(frac_Norm2[15]), .B(frac[18]), .C(n70739), 
         .D(n70613), .Z(n10673[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i16_4_lut.init = 16'hcac0;
    LUT4 i116_4_lut (.A(n8360[1]), .B(efectExp[1]), .C(n70739), .D(n40687), 
         .Z(n769)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i116_4_lut.init = 16'hcac0;
    LUT4 mux_52_i5_3_lut (.A(A_int[1]), .B(B_int[1]), .C(n70737), .Z(n480[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i5_3_lut.init = 16'hacac;
    LUT4 mux_51_i5_3_lut (.A(addSubAB[4]), .B(subBAExpEq[4]), .C(n70733), 
         .Z(n451[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i5_3_lut.init = 16'hcaca;
    LUT4 i55060_1_lut_4_lut (.A(n66206), .B(n9_c), .C(n14_adj_418), .D(n10_adj_419), 
         .Z(n67677)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i55060_1_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_rep_767 (.A(n66206), .B(n9_c), .C(n14_adj_418), .D(n10_adj_419), 
         .Z(n70737)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_rep_767.init = 16'hfffe;
    CCU2D sub_211_add_2_9 (.A0(B_int[30]), .B0(A_int[30]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61859), .S0(diffExpBA[7]), .S1(diffExpBA[8]));
    defparam sub_211_add_2_9.INIT0 = 16'h5999;
    defparam sub_211_add_2_9.INIT1 = 16'hffff;
    defparam sub_211_add_2_9.INJECT1_0 = "NO";
    defparam sub_211_add_2_9.INJECT1_1 = "NO";
    CCU2D equal_48_8 (.A0(B_int[24]), .B0(A_int[24]), .C0(B_int[23]), 
          .D0(A_int[23]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n60992), .S1(n448));
    defparam equal_48_8.INIT0 = 16'h9009;
    defparam equal_48_8.INIT1 = 16'hFFFF;
    defparam equal_48_8.INJECT1_0 = "YES";
    defparam equal_48_8.INJECT1_1 = "NO";
    LUT4 mux_52_i6_3_lut (.A(\A_int[2] ), .B(\B_int[2] ), .C(n70737), 
         .Z(n480[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i6_3_lut.init = 16'hacac;
    LUT4 i5_2_lut (.A(B_int[5]), .B(\B_int[3] ), .Z(n28_c)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    CCU2D sub_211_add_2_7 (.A0(B_int[28]), .B0(A_int[28]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[29]), .B1(A_int[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61858), .COUT(n61859), .S0(diffExpBA[5]), 
          .S1(diffExpBA[6]));
    defparam sub_211_add_2_7.INIT0 = 16'h5999;
    defparam sub_211_add_2_7.INIT1 = 16'h5999;
    defparam sub_211_add_2_7.INJECT1_0 = "NO";
    defparam sub_211_add_2_7.INJECT1_1 = "NO";
    FD1P3AX A_int_i0_i31 (.D(alu_a[31]), .SP(n73804), .CK(clock), .Q(A_int[31]));
    defparam A_int_i0_i31.GSR = "DISABLED";
    LUT4 mux_51_i6_3_lut (.A(addSubAB[5]), .B(subBAExpEq[5]), .C(n70733), 
         .Z(n451[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i6_3_lut.init = 16'hcaca;
    LUT4 mux_52_i4_3_lut (.A(A_int[0]), .B(B_int[0]), .C(n70737), .Z(n480[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i4_3_lut.init = 16'hacac;
    LUT4 mux_51_i4_3_lut (.A(addSubAB[3]), .B(subBAExpEq[3]), .C(n70733), 
         .Z(n451[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i4_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut (.A(frac[8]), .B(n70715), .C(frac[17]), .D(frac[23]), 
         .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(n31), .B(frac[18]), .C(n24), .D(n70805), .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(frac[24]), .B(frac[10]), .Z(n29)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i6_2_lut (.A(frac[9]), .B(frac[7]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i14_4_lut (.A(frac[11]), .B(frac[19]), .C(n70714), .D(n70703), 
         .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(n29), .B(n36), .C(n66182), .D(frac[6]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n41758)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    CCU2D sub_211_add_2_5 (.A0(B_int[26]), .B0(A_int[26]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[27]), .B1(A_int[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61857), .COUT(n61858), .S0(diffExpBA[3]), 
          .S1(diffExpBA[4]));
    defparam sub_211_add_2_5.INIT0 = 16'h5999;
    defparam sub_211_add_2_5.INIT1 = 16'h5999;
    defparam sub_211_add_2_5.INJECT1_0 = "NO";
    defparam sub_211_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_211_add_2_3 (.A0(B_int[24]), .B0(A_int[24]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[25]), .B1(A_int[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61856), .COUT(n61857), .S0(diffExpBA[1]), 
          .S1(diffExpBA[2]));
    defparam sub_211_add_2_3.INIT0 = 16'h5999;
    defparam sub_211_add_2_3.INIT1 = 16'h5999;
    defparam sub_211_add_2_3.INJECT1_0 = "NO";
    defparam sub_211_add_2_3.INJECT1_1 = "NO";
    FD1P3AX A_int_i0_i30 (.D(alu_a[30]), .SP(n73804), .CK(clock), .Q(A_int[30]));
    defparam A_int_i0_i30.GSR = "DISABLED";
    FD1P3AX A_int_i0_i29 (.D(alu_a[29]), .SP(n73804), .CK(clock), .Q(A_int[29]));
    defparam A_int_i0_i29.GSR = "DISABLED";
    FD1P3AX A_int_i0_i28 (.D(alu_a[28]), .SP(n73804), .CK(clock), .Q(A_int[28]));
    defparam A_int_i0_i28.GSR = "DISABLED";
    FD1P3AX A_int_i0_i27 (.D(alu_a[27]), .SP(n73804), .CK(clock), .Q(A_int[27]));
    defparam A_int_i0_i27.GSR = "DISABLED";
    FD1P3AX A_int_i0_i26 (.D(alu_a[26]), .SP(n73804), .CK(clock), .Q(A_int[26]));
    defparam A_int_i0_i26.GSR = "DISABLED";
    FD1P3AX A_int_i0_i25 (.D(alu_a[25]), .SP(n73804), .CK(clock), .Q(A_int[25]));
    defparam A_int_i0_i25.GSR = "DISABLED";
    FD1P3AX A_int_i0_i24 (.D(alu_a[24]), .SP(n73804), .CK(clock), .Q(A_int[24]));
    defparam A_int_i0_i24.GSR = "DISABLED";
    FD1P3AX A_int_i0_i23 (.D(alu_a[23]), .SP(n73804), .CK(clock), .Q(A_int[23]));
    defparam A_int_i0_i23.GSR = "DISABLED";
    FD1P3AX A_int_i0_i22 (.D(alu_a[22]), .SP(n73804), .CK(clock), .Q(A_int[22]));
    defparam A_int_i0_i22.GSR = "DISABLED";
    FD1P3AX A_int_i0_i21 (.D(alu_a[21]), .SP(n73804), .CK(clock), .Q(A_int[21]));
    defparam A_int_i0_i21.GSR = "DISABLED";
    FD1P3AX A_int_i0_i20 (.D(alu_a[20]), .SP(n73804), .CK(clock), .Q(A_int[20]));
    defparam A_int_i0_i20.GSR = "DISABLED";
    FD1P3AX A_int_i0_i19 (.D(alu_a[19]), .SP(n73804), .CK(clock), .Q(A_int[19]));
    defparam A_int_i0_i19.GSR = "DISABLED";
    FD1P3AX A_int_i0_i18 (.D(alu_a[18]), .SP(n73804), .CK(clock), .Q(\A_int[18] ));
    defparam A_int_i0_i18.GSR = "DISABLED";
    FD1P3AX A_int_i0_i17 (.D(alu_a[17]), .SP(n73804), .CK(clock), .Q(\A_int[17] ));
    defparam A_int_i0_i17.GSR = "DISABLED";
    FD1P3AX A_int_i0_i16 (.D(alu_a[16]), .SP(n73804), .CK(clock), .Q(\A_int[16] ));
    defparam A_int_i0_i16.GSR = "DISABLED";
    FD1P3AX A_int_i0_i15 (.D(alu_a[15]), .SP(n73804), .CK(clock), .Q(A_int[15]));
    defparam A_int_i0_i15.GSR = "DISABLED";
    FD1P3AX A_int_i0_i14 (.D(alu_a[14]), .SP(n73804), .CK(clock), .Q(A_int[14]));
    defparam A_int_i0_i14.GSR = "DISABLED";
    FD1P3AX A_int_i0_i13 (.D(alu_a[13]), .SP(n73804), .CK(clock), .Q(\A_int[13] ));
    defparam A_int_i0_i13.GSR = "DISABLED";
    FD1P3AX A_int_i0_i12 (.D(alu_a[12]), .SP(n73804), .CK(clock), .Q(\A_int[12] ));
    defparam A_int_i0_i12.GSR = "DISABLED";
    FD1P3AX A_int_i0_i11 (.D(alu_a[11]), .SP(n73804), .CK(clock), .Q(\A_int[11] ));
    defparam A_int_i0_i11.GSR = "DISABLED";
    FD1P3AX A_int_i0_i10 (.D(alu_a[10]), .SP(n73804), .CK(clock), .Q(\A_int[10] ));
    defparam A_int_i0_i10.GSR = "DISABLED";
    FD1P3AX A_int_i0_i9 (.D(alu_a[9]), .SP(n73804), .CK(clock), .Q(\A_int[9] ));
    defparam A_int_i0_i9.GSR = "DISABLED";
    FD1P3AX A_int_i0_i8 (.D(alu_a[8]), .SP(n73804), .CK(clock), .Q(A_int[8]));
    defparam A_int_i0_i8.GSR = "DISABLED";
    FD1P3AX A_int_i0_i7 (.D(alu_a[7]), .SP(n73804), .CK(clock), .Q(\A_int[7] ));
    defparam A_int_i0_i7.GSR = "DISABLED";
    FD1P3AX A_int_i0_i6 (.D(alu_a[6]), .SP(n73804), .CK(clock), .Q(A_int[6]));
    defparam A_int_i0_i6.GSR = "DISABLED";
    FD1P3AX A_int_i0_i5 (.D(alu_a[5]), .SP(n73804), .CK(clock), .Q(A_int[5]));
    defparam A_int_i0_i5.GSR = "DISABLED";
    FD1P3AX A_int_i0_i4 (.D(alu_a[4]), .SP(n73804), .CK(clock), .Q(\A_int[4] ));
    defparam A_int_i0_i4.GSR = "DISABLED";
    FD1P3AX A_int_i0_i3 (.D(alu_a[3]), .SP(n73804), .CK(clock), .Q(\A_int[3] ));
    defparam A_int_i0_i3.GSR = "DISABLED";
    FD1P3AX A_int_i0_i2 (.D(alu_a[2]), .SP(n73804), .CK(clock), .Q(\A_int[2] ));
    defparam A_int_i0_i2.GSR = "DISABLED";
    FD1P3AX A_int_i0_i1 (.D(alu_a[1]), .SP(n73804), .CK(clock), .Q(A_int[1]));
    defparam A_int_i0_i1.GSR = "DISABLED";
    FD1P3AX FP_Z_i0_i31 (.D(sign), .SP(n73804), .CK(clock), .Q(add_c[31]));
    defparam FP_Z_i0_i31.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_756_4_lut (.A(n70805), .B(subBAExpEq[27]), .C(n448), 
         .D(n70739), .Z(n70726)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_2_lut_rep_756_4_lut.init = 16'hff10;
    FD1P3AX B_int_i0_i31 (.D(alu_b[31]), .SP(add_ce), .CK(clock), .Q(B_int[31]));
    defparam B_int_i0_i31.GSR = "DISABLED";
    FD1P3AX B_int_i0_i30 (.D(alu_b[30]), .SP(add_ce), .CK(clock), .Q(B_int[30]));
    defparam B_int_i0_i30.GSR = "DISABLED";
    FD1P3AX B_int_i0_i29 (.D(alu_b[29]), .SP(add_ce), .CK(clock), .Q(B_int[29]));
    defparam B_int_i0_i29.GSR = "DISABLED";
    FD1P3AX B_int_i0_i28 (.D(alu_b[28]), .SP(add_ce), .CK(clock), .Q(B_int[28]));
    defparam B_int_i0_i28.GSR = "DISABLED";
    FD1P3AX B_int_i0_i27 (.D(alu_b[27]), .SP(add_ce), .CK(clock), .Q(B_int[27]));
    defparam B_int_i0_i27.GSR = "DISABLED";
    FD1P3AX B_int_i0_i26 (.D(alu_b[26]), .SP(add_ce), .CK(clock), .Q(B_int[26]));
    defparam B_int_i0_i26.GSR = "DISABLED";
    FD1P3AX B_int_i0_i25 (.D(alu_b[25]), .SP(add_ce), .CK(clock), .Q(B_int[25]));
    defparam B_int_i0_i25.GSR = "DISABLED";
    FD1P3AX B_int_i0_i24 (.D(alu_b[24]), .SP(add_ce), .CK(clock), .Q(B_int[24]));
    defparam B_int_i0_i24.GSR = "DISABLED";
    FD1P3AX B_int_i0_i23 (.D(alu_b[23]), .SP(add_ce), .CK(clock), .Q(B_int[23]));
    defparam B_int_i0_i23.GSR = "DISABLED";
    FD1P3AX B_int_i0_i22 (.D(alu_b[22]), .SP(add_ce), .CK(clock), .Q(B_int[22]));
    defparam B_int_i0_i22.GSR = "DISABLED";
    FD1P3AX B_int_i0_i21 (.D(alu_b[21]), .SP(add_ce), .CK(clock), .Q(B_int[21]));
    defparam B_int_i0_i21.GSR = "DISABLED";
    FD1P3AX B_int_i0_i20 (.D(alu_b[20]), .SP(add_ce), .CK(clock), .Q(B_int[20]));
    defparam B_int_i0_i20.GSR = "DISABLED";
    FD1P3AX B_int_i0_i19 (.D(alu_b[19]), .SP(add_ce), .CK(clock), .Q(B_int[19]));
    defparam B_int_i0_i19.GSR = "DISABLED";
    FD1P3AX B_int_i0_i18 (.D(alu_b[18]), .SP(add_ce), .CK(clock), .Q(\B_int[18] ));
    defparam B_int_i0_i18.GSR = "DISABLED";
    FD1P3AX B_int_i0_i17 (.D(alu_b[17]), .SP(add_ce), .CK(clock), .Q(\B_int[17] ));
    defparam B_int_i0_i17.GSR = "DISABLED";
    FD1P3AX B_int_i0_i16 (.D(alu_b[16]), .SP(add_ce), .CK(clock), .Q(\B_int[16] ));
    defparam B_int_i0_i16.GSR = "DISABLED";
    FD1P3AX B_int_i0_i15 (.D(alu_b[15]), .SP(add_ce), .CK(clock), .Q(B_int[15]));
    defparam B_int_i0_i15.GSR = "DISABLED";
    FD1P3AX B_int_i0_i14 (.D(alu_b[14]), .SP(add_ce), .CK(clock), .Q(B_int[14]));
    defparam B_int_i0_i14.GSR = "DISABLED";
    FD1P3AX B_int_i0_i13 (.D(alu_b[13]), .SP(add_ce), .CK(clock), .Q(\B_int[13] ));
    defparam B_int_i0_i13.GSR = "DISABLED";
    FD1P3AX B_int_i0_i12 (.D(alu_b[12]), .SP(add_ce), .CK(clock), .Q(\B_int[12] ));
    defparam B_int_i0_i12.GSR = "DISABLED";
    FD1P3AX B_int_i0_i11 (.D(alu_b[11]), .SP(add_ce), .CK(clock), .Q(\B_int[11] ));
    defparam B_int_i0_i11.GSR = "DISABLED";
    FD1P3AX B_int_i0_i10 (.D(alu_b[10]), .SP(add_ce), .CK(clock), .Q(\B_int[10] ));
    defparam B_int_i0_i10.GSR = "DISABLED";
    FD1P3AX B_int_i0_i9 (.D(alu_b[9]), .SP(add_ce), .CK(clock), .Q(\B_int[9] ));
    defparam B_int_i0_i9.GSR = "DISABLED";
    FD1P3AX B_int_i0_i8 (.D(alu_b[8]), .SP(add_ce), .CK(clock), .Q(B_int[8]));
    defparam B_int_i0_i8.GSR = "DISABLED";
    FD1P3AX B_int_i0_i7 (.D(alu_b[7]), .SP(add_ce), .CK(clock), .Q(\B_int[7] ));
    defparam B_int_i0_i7.GSR = "DISABLED";
    FD1P3AX B_int_i0_i6 (.D(alu_b[6]), .SP(add_ce), .CK(clock), .Q(B_int[6]));
    defparam B_int_i0_i6.GSR = "DISABLED";
    FD1P3AX B_int_i0_i5 (.D(alu_b[5]), .SP(add_ce), .CK(clock), .Q(B_int[5]));
    defparam B_int_i0_i5.GSR = "DISABLED";
    FD1P3AX B_int_i0_i4 (.D(alu_b[4]), .SP(add_ce), .CK(clock), .Q(\B_int[4] ));
    defparam B_int_i0_i4.GSR = "DISABLED";
    FD1P3AX B_int_i0_i3 (.D(alu_b[3]), .SP(add_ce), .CK(clock), .Q(\B_int[3] ));
    defparam B_int_i0_i3.GSR = "DISABLED";
    FD1P3AX B_int_i0_i2 (.D(alu_b[2]), .SP(add_ce), .CK(clock), .Q(\B_int[2] ));
    defparam B_int_i0_i2.GSR = "DISABLED";
    FD1P3AX B_int_i0_i1 (.D(alu_b[1]), .SP(add_ce), .CK(clock), .Q(B_int[1]));
    defparam B_int_i0_i1.GSR = "DISABLED";
    LUT4 i117_4_lut (.A(n8360[0]), .B(efectExp[0]), .C(n70739), .D(n40687), 
         .Z(n770)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i117_4_lut.init = 16'hcac0;
    LUT4 i15_4_lut (.A(\B_int[7] ), .B(B_int[22]), .C(\B_int[4] ), .D(B_int[14]), 
         .Z(n38_adj_420)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 mux_3773_i4_4_lut (.A(frac_Norm2[3]), .B(frac[6]), .C(n70739), 
         .D(n70613), .Z(n10673[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i4_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i3_4_lut (.A(frac_Norm2[2]), .B(n70703), .C(n70739), 
         .D(n70613), .Z(n10673[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i3_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i2_4_lut (.A(frac_Norm2[1]), .B(n70706), .C(n70739), 
         .D(n70613), .Z(n10673[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i2_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut (.A(B_int[21]), .B(B_int[1]), .Z(n24_adj_421)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i13_4_lut (.A(\B_int[2] ), .B(B_int[20]), .C(\B_int[17] ), .D(\B_int[12] ), 
         .Z(n36_adj_422)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut_adj_781 (.A(B_int[0]), .B(n38_adj_420), .C(n28_c), 
         .D(\B_int[9] ), .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_781.init = 16'hfffe;
    LUT4 i9_2_lut_adj_782 (.A(\B_int[18] ), .B(\B_int[11] ), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut_adj_782.init = 16'heeee;
    CCU2D sub_211_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(B_int[23]), .B1(A_int[23]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61856), .S1(diffExpBA[0]));
    defparam sub_211_add_2_1.INIT0 = 16'h0000;
    defparam sub_211_add_2_1.INIT1 = 16'h5999;
    defparam sub_211_add_2_1.INJECT1_0 = "NO";
    defparam sub_211_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_668_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n39), 
         .D(n70643), .Z(n70638)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_668_4_lut_4_lut.init = 16'h8000;
    LUT4 mux_3773_i23_4_lut (.A(frac_Norm2[22]), .B(frac[25]), .C(n70739), 
         .D(n70613), .Z(n10673[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i23_4_lut.init = 16'hcac0;
    LUT4 i28246_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(frac[12]), 
         .D(n39), .Z(n243[12])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28246_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(\B_int[10] ), .B(B_int[15]), .C(B_int[6]), .D(B_int[19]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i29393_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n19140), 
         .D(n39), .Z(n272[10])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i29393_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    CCU2D equal_48_7 (.A0(B_int[28]), .B0(A_int[28]), .C0(B_int[27]), 
          .D0(A_int[27]), .A1(B_int[26]), .B1(A_int[26]), .C1(B_int[25]), 
          .D1(A_int[25]), .CIN(n60991), .COUT(n60992));
    defparam equal_48_7.INIT0 = 16'h9009;
    defparam equal_48_7.INIT1 = 16'h9009;
    defparam equal_48_7.INJECT1_0 = "YES";
    defparam equal_48_7.INJECT1_1 = "YES";
    LUT4 i1_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n70707), 
         .D(n39), .Z(n4)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    FD1P3IX FP_Z_i0_i1 (.D(n10673[1]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[1]));
    defparam FP_Z_i0_i1.GSR = "DISABLED";
    LUT4 i28250_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(frac[8]), 
         .D(n39), .Z(n243[8])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28250_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    FD1P3IX FP_Z_i0_i2 (.D(n10673[2]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[2]));
    defparam FP_Z_i0_i2.GSR = "DISABLED";
    LUT4 i28247_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(frac[11]), 
         .D(n39), .Z(n243[11])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28247_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 i21_4_lut (.A(\B_int[13] ), .B(n42), .C(n36_adj_422), .D(n24_adj_421), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    FD1P3IX FP_Z_i0_i3 (.D(n10673[3]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[3]));
    defparam FP_Z_i0_i3.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_666_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), 
         .C(efectExp[4]), .D(n39), .Z(n70636)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_rep_666_4_lut_4_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_rep_667_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), 
         .C(n70726), .D(n39), .Z(n70637)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_667_4_lut_4_lut_4_lut.init = 16'hf7ff;
    LUT4 i110_4_lut (.A(n8360[7]), .B(efectExp[7]), .C(n70739), .D(n40687), 
         .Z(n763)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i110_4_lut.init = 16'hcac0;
    LUT4 i111_4_lut (.A(n8360[6]), .B(efectExp[6]), .C(n70739), .D(n40687), 
         .Z(n764)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i111_4_lut.init = 16'hcac0;
    LUT4 i112_4_lut (.A(n8360[5]), .B(efectExp[5]), .C(n70739), .D(n40687), 
         .Z(n765)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i112_4_lut.init = 16'hcac0;
    LUT4 i28409_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n70805), 
         .D(n39), .Z(n40002)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i28409_2_lut_4_lut_4_lut_4_lut.init = 16'hf7ff;
    LUT4 i8_2_lut (.A(B_int[8]), .B(\B_int[16] ), .Z(n31_adj_424)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i22_4_lut (.A(n31_adj_424), .B(n44), .C(n40), .D(n32), .Z(n66192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut_adj_783 (.A(A_int[15]), .B(A_int[14]), .Z(n28_adj_425)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut_adj_783.init = 16'heeee;
    LUT4 i15_4_lut_adj_784 (.A(\A_int[16] ), .B(A_int[21]), .C(\A_int[3] ), 
         .D(\A_int[18] ), .Z(n38_adj_426)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut_adj_784.init = 16'hfffe;
    LUT4 i1_2_lut_adj_785 (.A(A_int[1]), .B(\A_int[12] ), .Z(n24_adj_427)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_785.init = 16'heeee;
    LUT4 i2_2_lut_adj_786 (.A(A_int[27]), .B(A_int[23]), .Z(n10_adj_428)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_786.init = 16'h8888;
    LUT4 i28245_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(frac[13]), 
         .D(n39), .Z(n243[13])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28245_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    CCU2D equal_48_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(B_int[30]), .B1(A_int[30]), .C1(B_int[29]), .D1(A_int[29]), 
          .COUT(n60991));
    defparam equal_48_0.INIT0 = 16'hF000;
    defparam equal_48_0.INIT1 = 16'h9009;
    defparam equal_48_0.INJECT1_0 = "NO";
    defparam equal_48_0.INJECT1_1 = "YES";
    LUT4 i28248_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(frac[10]), 
         .D(n39), .Z(n243[10])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28248_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 mux_3773_i19_4_lut (.A(frac_Norm2[18]), .B(frac[21]), .C(n70739), 
         .D(n70613), .Z(n10673[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i19_4_lut.init = 16'hcac0;
    LUT4 i113_4_lut (.A(n8360[4]), .B(efectExp[4]), .C(n70739), .D(n40687), 
         .Z(n766)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i113_4_lut.init = 16'hcac0;
    LUT4 mux_3773_i18_4_lut (.A(frac_Norm2[17]), .B(frac[20]), .C(n70739), 
         .D(n70613), .Z(n10673[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i18_4_lut.init = 16'hcac0;
    LUT4 i28251_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(frac[6]), 
         .D(n39), .Z(n243[6])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28251_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 i13_4_lut_adj_787 (.A(A_int[0]), .B(\A_int[10] ), .C(A_int[19]), 
         .D(A_int[6]), .Z(n36_adj_429)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_787.init = 16'hfffe;
    LUT4 i19_4_lut_adj_788 (.A(\A_int[4] ), .B(n38_adj_426), .C(n28_adj_425), 
         .D(A_int[22]), .Z(n42_adj_430)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_788.init = 16'hfffe;
    LUT4 i29394_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n19142), 
         .D(n39), .Z(n272[9])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i29394_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 i9_2_lut_adj_789 (.A(A_int[20]), .B(A_int[8]), .Z(n32_adj_431)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut_adj_789.init = 16'heeee;
    FD1P3IX FP_Z_i0_i4 (.D(n10673[4]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[4]));
    defparam FP_Z_i0_i4.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i5 (.D(n10673[5]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[5]));
    defparam FP_Z_i0_i5.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i6 (.D(n10673[6]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[6]));
    defparam FP_Z_i0_i6.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i7 (.D(n10673[7]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[7]));
    defparam FP_Z_i0_i7.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i8 (.D(n10673[8]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[8]));
    defparam FP_Z_i0_i8.GSR = "DISABLED";
    LUT4 i17_4_lut_adj_790 (.A(\A_int[17] ), .B(\A_int[2] ), .C(A_int[5]), 
         .D(\A_int[13] ), .Z(n40_adj_432)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_790.init = 16'hfffe;
    LUT4 i28252_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n70703), 
         .D(n39), .Z(n243[5])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28252_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 i21_4_lut_adj_791 (.A(\A_int[9] ), .B(n42_adj_430), .C(n36_adj_429), 
         .D(n24_adj_427), .Z(n44_adj_433)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut_adj_791.init = 16'hfffe;
    LUT4 i8_2_lut_adj_792 (.A(\A_int[11] ), .B(\A_int[7] ), .Z(n31_adj_434)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut_adj_792.init = 16'heeee;
    FD1P3IX FP_Z_i0_i9 (.D(n10673[9]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[9]));
    defparam FP_Z_i0_i9.GSR = "DISABLED";
    LUT4 i22_4_lut_adj_793 (.A(n31_adj_434), .B(n44_adj_433), .C(n40_adj_432), 
         .D(n32_adj_431), .Z(n66206)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut_adj_793.init = 16'hfffe;
    FD1P3IX FP_Z_i0_i10 (.D(n10673[10]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[10]));
    defparam FP_Z_i0_i10.GSR = "DISABLED";
    LUT4 i2_2_lut_adj_794 (.A(A_int[24]), .B(A_int[30]), .Z(n10_adj_419)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_794.init = 16'heeee;
    LUT4 i6_4_lut_adj_795 (.A(A_int[28]), .B(A_int[23]), .C(A_int[26]), 
         .D(A_int[27]), .Z(n14_adj_418)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_795.init = 16'hfffe;
    LUT4 i1_2_lut_adj_796 (.A(A_int[25]), .B(A_int[29]), .Z(n9_c)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_796.init = 16'heeee;
    LUT4 i29392_2_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n19138), 
         .D(n39), .Z(n272[11])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i29392_2_lut_4_lut_4_lut_4_lut.init = 16'h8000;
    LUT4 i8759_2_lut_rep_663_4_lut_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), 
         .C(n66653), .D(n39), .Z(n70633)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i8759_2_lut_rep_663_4_lut_4_lut_4_lut_4_lut.init = 16'h7fff;
    FD1P3IX FP_Z_i0_i11 (.D(n10673[11]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[11]));
    defparam FP_Z_i0_i11.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i12 (.D(n10673[12]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[12]));
    defparam FP_Z_i0_i12.GSR = "DISABLED";
    LUT4 i6_4_lut_adj_797 (.A(A_int[26]), .B(A_int[25]), .C(A_int[28]), 
         .D(A_int[30]), .Z(n14_adj_435)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_797.init = 16'h8000;
    FD1P3IX FP_Z_i0_i13 (.D(n10673[13]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[13]));
    defparam FP_Z_i0_i13.GSR = "DISABLED";
    FD1P3IX FP_Z_i0_i14 (.D(n10673[14]), .SP(add_ce), .CD(n24122), .CK(clock), 
            .Q(add_c[14]));
    defparam FP_Z_i0_i14.GSR = "DISABLED";
    LUT4 i1_4_lut_rep_899_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n66653), 
         .D(n39), .Z(n73795)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;
    defparam i1_4_lut_rep_899_4_lut_4_lut.init = 16'h3b33;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n31_adj_423), .B(n70641), .C(n21808), 
         .D(n39), .Z(leadZerosBin[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A !((D)+!B)) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'h80cc;
    PFUMX i29 (.BLUT(n66558), .ALUT(n19), .C0(isSUB), .Z(n63661));
    PFUMX i28 (.BLUT(n15), .ALUT(n18), .C0(isSUB), .Z(n63665));
    PFUMX mux_215_i3 (.BLUT(frac_add_Norm1[2]), .ALUT(frac_sub_Norm1[2]), 
          .C0(isSUB), .Z(frac_Norm1[2]));
    PFUMX mux_215_i4 (.BLUT(frac_add_Norm1[3]), .ALUT(frac_sub_Norm1[3]), 
          .C0(isSUB), .Z(frac_Norm1[3]));
    CCU2D sub_214_add_2_25 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61531), .S0(subBAExpEq[26]), .S1(subBAExpEq[27]));
    defparam sub_214_add_2_25.INIT0 = 16'h0fff;
    defparam sub_214_add_2_25.INIT1 = 16'hffff;
    defparam sub_214_add_2_25.INJECT1_0 = "NO";
    defparam sub_214_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_23 (.A0(B_int[21]), .B0(A_int[21]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[22]), .B1(A_int[22]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61530), .COUT(n61531), .S0(subBAExpEq[24]), 
          .S1(subBAExpEq[25]));
    defparam sub_214_add_2_23.INIT0 = 16'h5999;
    defparam sub_214_add_2_23.INIT1 = 16'h5999;
    defparam sub_214_add_2_23.INJECT1_0 = "NO";
    defparam sub_214_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_21 (.A0(B_int[19]), .B0(A_int[19]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[20]), .B1(A_int[20]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61529), .COUT(n61530), .S0(subBAExpEq[22]), 
          .S1(subBAExpEq[23]));
    defparam sub_214_add_2_21.INIT0 = 16'h5999;
    defparam sub_214_add_2_21.INIT1 = 16'h5999;
    defparam sub_214_add_2_21.INJECT1_0 = "NO";
    defparam sub_214_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_19 (.A0(\B_int[17] ), .B0(\A_int[17] ), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[18] ), .B1(\A_int[18] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61528), .COUT(n61529), .S0(subBAExpEq[20]), 
          .S1(subBAExpEq[21]));
    defparam sub_214_add_2_19.INIT0 = 16'h5999;
    defparam sub_214_add_2_19.INIT1 = 16'h5999;
    defparam sub_214_add_2_19.INJECT1_0 = "NO";
    defparam sub_214_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_17 (.A0(B_int[15]), .B0(A_int[15]), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[16] ), .B1(\A_int[16] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61527), .COUT(n61528), .S0(subBAExpEq[18]), 
          .S1(subBAExpEq[19]));
    defparam sub_214_add_2_17.INIT0 = 16'h5999;
    defparam sub_214_add_2_17.INIT1 = 16'h5999;
    defparam sub_214_add_2_17.INJECT1_0 = "NO";
    defparam sub_214_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_15 (.A0(\B_int[13] ), .B0(\A_int[13] ), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[14]), .B1(A_int[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61526), .COUT(n61527), .S0(subBAExpEq[16]), 
          .S1(subBAExpEq[17]));
    defparam sub_214_add_2_15.INIT0 = 16'h5999;
    defparam sub_214_add_2_15.INIT1 = 16'h5999;
    defparam sub_214_add_2_15.INJECT1_0 = "NO";
    defparam sub_214_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_13 (.A0(\B_int[11] ), .B0(\A_int[11] ), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[12] ), .B1(\A_int[12] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61525), .COUT(n61526), .S0(subBAExpEq[14]), 
          .S1(subBAExpEq[15]));
    defparam sub_214_add_2_13.INIT0 = 16'h5999;
    defparam sub_214_add_2_13.INIT1 = 16'h5999;
    defparam sub_214_add_2_13.INJECT1_0 = "NO";
    defparam sub_214_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_11 (.A0(\B_int[9] ), .B0(\A_int[9] ), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[10] ), .B1(\A_int[10] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61524), .COUT(n61525), .S0(subBAExpEq[12]), 
          .S1(subBAExpEq[13]));
    defparam sub_214_add_2_11.INIT0 = 16'h5999;
    defparam sub_214_add_2_11.INIT1 = 16'h5999;
    defparam sub_214_add_2_11.INJECT1_0 = "NO";
    defparam sub_214_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_9 (.A0(\B_int[7] ), .B0(\A_int[7] ), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[8]), .B1(A_int[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61523), .COUT(n61524), .S0(subBAExpEq[10]), 
          .S1(subBAExpEq[11]));
    defparam sub_214_add_2_9.INIT0 = 16'h5999;
    defparam sub_214_add_2_9.INIT1 = 16'h5999;
    defparam sub_214_add_2_9.INJECT1_0 = "NO";
    defparam sub_214_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_7 (.A0(B_int[5]), .B0(A_int[5]), .C0(GND_net), 
          .D0(GND_net), .A1(B_int[6]), .B1(A_int[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61522), .COUT(n61523), .S0(subBAExpEq[8]), 
          .S1(subBAExpEq[9]));
    defparam sub_214_add_2_7.INIT0 = 16'h5999;
    defparam sub_214_add_2_7.INIT1 = 16'h5999;
    defparam sub_214_add_2_7.INJECT1_0 = "NO";
    defparam sub_214_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_5 (.A0(\B_int[3] ), .B0(\A_int[3] ), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[4] ), .B1(\A_int[4] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61521), .COUT(n61522), .S0(subBAExpEq[6]), 
          .S1(subBAExpEq[7]));
    defparam sub_214_add_2_5.INIT0 = 16'h5999;
    defparam sub_214_add_2_5.INIT1 = 16'h5999;
    defparam sub_214_add_2_5.INJECT1_0 = "NO";
    defparam sub_214_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_214_add_2_3 (.A0(B_int[1]), .B0(A_int[1]), .C0(GND_net), 
          .D0(GND_net), .A1(\B_int[2] ), .B1(\A_int[2] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n61520), .COUT(n61521), .S0(subBAExpEq[4]), 
          .S1(subBAExpEq[5]));
    defparam sub_214_add_2_3.INIT0 = 16'h5999;
    defparam sub_214_add_2_3.INIT1 = 16'h5999;
    defparam sub_214_add_2_3.INJECT1_0 = "NO";
    defparam sub_214_add_2_3.INJECT1_1 = "NO";
    LUT4 i6694_2_lut (.A(addSubAB[27]), .B(diffExpAB[8]), .Z(n17318)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6694_2_lut.init = 16'heeee;
    CCU2D sub_214_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(B_int[0]), .B1(A_int[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61520), .S1(subBAExpEq[3]));
    defparam sub_214_add_2_1.INIT0 = 16'h0000;
    defparam sub_214_add_2_1.INIT1 = 16'h5999;
    defparam sub_214_add_2_1.INJECT1_0 = "NO";
    defparam sub_214_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_9 (.A0(A_int[30]), .B0(B_int[30]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61518), .S0(diffExpAB_c[7]), .S1(diffExpAB[8]));
    defparam sub_210_add_2_9.INIT0 = 16'h5999;
    defparam sub_210_add_2_9.INIT1 = 16'hffff;
    defparam sub_210_add_2_9.INJECT1_0 = "NO";
    defparam sub_210_add_2_9.INJECT1_1 = "NO";
    CCU2D add_3092_29 (.A0(A_int[31]), .B0(n70865), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62218), 
          .S0(addSubAB[27]));
    defparam add_3092_29.INIT0 = 16'h6999;
    defparam add_3092_29.INIT1 = 16'h0000;
    defparam add_3092_29.INJECT1_0 = "NO";
    defparam add_3092_29.INJECT1_1 = "NO";
    CCU2D add_3092_27 (.A0(n21643), .B0(A_int[22]), .C0(B_int[22]), .D0(diffExpAB[8]), 
          .A1(n70805), .B1(n66178), .C1(GND_net), .D1(GND_net), .CIN(n62217), 
          .COUT(n62218), .S0(addSubAB[25]), .S1(addSubAB[26]));
    defparam add_3092_27.INIT0 = 16'ha599;
    defparam add_3092_27.INIT1 = 16'h9999;
    defparam add_3092_27.INJECT1_0 = "NO";
    defparam add_3092_27.INJECT1_1 = "NO";
    CCU2D add_3092_25 (.A0(n21651), .B0(A_int[20]), .C0(B_int[20]), .D0(diffExpAB[8]), 
          .A1(n21645), .B1(A_int[21]), .C1(B_int[21]), .D1(diffExpAB[8]), 
          .CIN(n62216), .COUT(n62217), .S0(addSubAB[23]), .S1(addSubAB[24]));
    defparam add_3092_25.INIT0 = 16'ha599;
    defparam add_3092_25.INIT1 = 16'ha599;
    defparam add_3092_25.INJECT1_0 = "NO";
    defparam add_3092_25.INJECT1_1 = "NO";
    LUT4 i6_4_lut_adj_798 (.A(B_int[23]), .B(B_int[24]), .C(B_int[27]), 
         .D(B_int[28]), .Z(n14_adj_436)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_798.init = 16'hfffe;
    LUT4 i5_4_lut (.A(B_int[25]), .B(B_int[29]), .C(B_int[30]), .D(B_int[26]), 
         .Z(n13)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    CCU2D add_3092_23 (.A0(n21681), .B0(\A_int[18] ), .C0(diffExpAB[8]), 
          .D0(\B_int[18] ), .A1(n21641), .B1(A_int[19]), .C1(B_int[19]), 
          .D1(diffExpAB[8]), .CIN(n62215), .COUT(n62216), .S0(addSubAB[21]), 
          .S1(addSubAB[22]));
    defparam add_3092_23.INIT0 = 16'ha959;
    defparam add_3092_23.INIT1 = 16'ha599;
    defparam add_3092_23.INJECT1_0 = "NO";
    defparam add_3092_23.INJECT1_1 = "NO";
    CCU2D add_3092_21 (.A0(n21679), .B0(diffExpAB[8]), .C0(\A_int[16] ), 
          .D0(\B_int[16] ), .A1(n21647), .B1(diffExpAB[8]), .C1(\B_int[17] ), 
          .D1(\A_int[17] ), .CIN(n62214), .COUT(n62215), .S0(addSubAB[19]), 
          .S1(addSubAB[20]));
    defparam add_3092_21.INIT0 = 16'ha965;
    defparam add_3092_21.INIT1 = 16'ha695;
    defparam add_3092_21.INJECT1_0 = "NO";
    defparam add_3092_21.INJECT1_1 = "NO";
    CCU2D add_3092_19 (.A0(n21665), .B0(A_int[14]), .C0(B_int[14]), .D0(diffExpAB[8]), 
          .A1(n21655), .B1(A_int[15]), .C1(B_int[15]), .D1(diffExpAB[8]), 
          .CIN(n62213), .COUT(n62214), .S0(addSubAB[17]), .S1(addSubAB[18]));
    defparam add_3092_19.INIT0 = 16'ha599;
    defparam add_3092_19.INIT1 = 16'ha599;
    defparam add_3092_19.INJECT1_0 = "NO";
    defparam add_3092_19.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_7 (.A0(A_int[28]), .B0(B_int[28]), .C0(GND_net), 
          .D0(GND_net), .A1(A_int[29]), .B1(B_int[29]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61517), .COUT(n61518), .S0(diffExpAB_c[5]), 
          .S1(diffExpAB_c[6]));
    defparam sub_210_add_2_7.INIT0 = 16'h5999;
    defparam sub_210_add_2_7.INIT1 = 16'h5999;
    defparam sub_210_add_2_7.INJECT1_0 = "NO";
    defparam sub_210_add_2_7.INJECT1_1 = "NO";
    CCU2D add_3092_17 (.A0(n21653), .B0(diffExpAB[8]), .C0(\B_int[12] ), 
          .D0(\A_int[12] ), .A1(n21667), .B1(diffExpAB[8]), .C1(\B_int[13] ), 
          .D1(\A_int[13] ), .CIN(n62212), .COUT(n62213), .S0(addSubAB[15]), 
          .S1(addSubAB[16]));
    defparam add_3092_17.INIT0 = 16'ha695;
    defparam add_3092_17.INIT1 = 16'ha695;
    defparam add_3092_17.INJECT1_0 = "NO";
    defparam add_3092_17.INJECT1_1 = "NO";
    CCU2D add_3092_15 (.A0(n21671), .B0(\A_int[10] ), .C0(diffExpAB[8]), 
          .D0(\B_int[10] ), .A1(n21657), .B1(diffExpAB[8]), .C1(\B_int[11] ), 
          .D1(\A_int[11] ), .CIN(n62211), .COUT(n62212), .S0(addSubAB[13]), 
          .S1(addSubAB[14]));
    defparam add_3092_15.INIT0 = 16'ha959;
    defparam add_3092_15.INIT1 = 16'ha695;
    defparam add_3092_15.INJECT1_0 = "NO";
    defparam add_3092_15.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_5 (.A0(A_int[26]), .B0(B_int[26]), .C0(GND_net), 
          .D0(GND_net), .A1(A_int[27]), .B1(B_int[27]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61516), .COUT(n61517), .S0(diffExpAB_c[3]), 
          .S1(diffExpAB_c[4]));
    defparam sub_210_add_2_5.INIT0 = 16'h5999;
    defparam sub_210_add_2_5.INIT1 = 16'h5999;
    defparam sub_210_add_2_5.INJECT1_0 = "NO";
    defparam sub_210_add_2_5.INJECT1_1 = "NO";
    CCU2D add_3092_13 (.A0(n21669), .B0(A_int[8]), .C0(B_int[8]), .D0(diffExpAB[8]), 
          .A1(n21677), .B1(diffExpAB[8]), .C1(\B_int[9] ), .D1(\A_int[9] ), 
          .CIN(n62210), .COUT(n62211), .S0(addSubAB[11]), .S1(addSubAB[12]));
    defparam add_3092_13.INIT0 = 16'ha599;
    defparam add_3092_13.INIT1 = 16'ha695;
    defparam add_3092_13.INJECT1_0 = "NO";
    defparam add_3092_13.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_3 (.A0(A_int[24]), .B0(B_int[24]), .C0(GND_net), 
          .D0(GND_net), .A1(A_int[25]), .B1(B_int[25]), .C1(GND_net), 
          .D1(GND_net), .CIN(n61515), .COUT(n61516), .S0(diffExpAB_c[1]), 
          .S1(diffExpAB_c[2]));
    defparam sub_210_add_2_3.INIT0 = 16'h5999;
    defparam sub_210_add_2_3.INIT1 = 16'h5999;
    defparam sub_210_add_2_3.INJECT1_0 = "NO";
    defparam sub_210_add_2_3.INJECT1_1 = "NO";
    CCU2D add_3092_11 (.A0(n21659), .B0(A_int[6]), .C0(B_int[6]), .D0(diffExpAB[8]), 
          .A1(n21663), .B1(diffExpAB[8]), .C1(\B_int[7] ), .D1(\A_int[7] ), 
          .CIN(n62209), .COUT(n62210), .S0(addSubAB[9]), .S1(addSubAB[10]));
    defparam add_3092_11.INIT0 = 16'ha599;
    defparam add_3092_11.INIT1 = 16'ha695;
    defparam add_3092_11.INJECT1_0 = "NO";
    defparam add_3092_11.INJECT1_1 = "NO";
    CCU2D add_3092_9 (.A0(n21661), .B0(\A_int[4] ), .C0(diffExpAB[8]), 
          .D0(\B_int[4] ), .A1(n21675), .B1(A_int[5]), .C1(B_int[5]), 
          .D1(diffExpAB[8]), .CIN(n62208), .COUT(n62209), .S0(addSubAB[7]), 
          .S1(addSubAB[8]));
    defparam add_3092_9.INIT0 = 16'ha959;
    defparam add_3092_9.INIT1 = 16'ha599;
    defparam add_3092_9.INJECT1_0 = "NO";
    defparam add_3092_9.INJECT1_1 = "NO";
    CCU2D add_3092_7 (.A0(n21687), .B0(diffExpAB[8]), .C0(\B_int[2] ), 
          .D0(\A_int[2] ), .A1(n21685), .B1(diffExpAB[8]), .C1(\B_int[3] ), 
          .D1(\A_int[3] ), .CIN(n62207), .COUT(n62208), .S0(addSubAB[5]), 
          .S1(addSubAB[6]));
    defparam add_3092_7.INIT0 = 16'ha695;
    defparam add_3092_7.INIT1 = 16'ha695;
    defparam add_3092_7.INJECT1_0 = "NO";
    defparam add_3092_7.INJECT1_1 = "NO";
    CCU2D add_3092_5 (.A0(n21711), .B0(A_int[0]), .C0(B_int[0]), .D0(diffExpAB[8]), 
          .A1(n21713), .B1(A_int[1]), .C1(B_int[1]), .D1(diffExpAB[8]), 
          .CIN(n62206), .COUT(n62207), .S0(addSubAB[3]), .S1(addSubAB[4]));
    defparam add_3092_5.INIT0 = 16'ha599;
    defparam add_3092_5.INIT1 = 16'ha599;
    defparam add_3092_5.INJECT1_0 = "NO";
    defparam add_3092_5.INJECT1_1 = "NO";
    LUT4 i7_4_lut_adj_799 (.A(A_int[24]), .B(n14_adj_435), .C(n10_adj_428), 
         .D(A_int[29]), .Z(expA_FF)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_799.init = 16'h8000;
    CCU2D add_3092_3 (.A0(efectFracB_align[1]), .B0(n70805), .C0(GND_net), 
          .D0(GND_net), .A1(efectFracB_align[2]), .B1(n70805), .C1(GND_net), 
          .D1(GND_net), .CIN(n62205), .COUT(n62206), .S0(addSubAB[1]), 
          .S1(addSubAB[2]));
    defparam add_3092_3.INIT0 = 16'h6999;
    defparam add_3092_3.INIT1 = 16'h6999;
    defparam add_3092_3.INJECT1_0 = "NO";
    defparam add_3092_3.INJECT1_1 = "NO";
    CCU2D add_3092_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(isSUB), .B1(n7), .C1(fracAlign_int[0]), .D1(n70805), .COUT(n62205), 
          .S1(addSubAB[0]));
    defparam add_3092_1.INIT0 = 16'hF000;
    defparam add_3092_1.INIT1 = 16'h56a9;
    defparam add_3092_1.INJECT1_0 = "NO";
    defparam add_3092_1.INJECT1_1 = "NO";
    CCU2D sub_210_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[23]), .B1(B_int[23]), .C1(GND_net), .D1(GND_net), 
          .COUT(n61515), .S1(diffExpAB_c[0]));
    defparam sub_210_add_2_1.INIT0 = 16'h0000;
    defparam sub_210_add_2_1.INIT1 = 16'h5999;
    defparam sub_210_add_2_1.INJECT1_0 = "NO";
    defparam sub_210_add_2_1.INJECT1_1 = "NO";
    CCU2D add_72_23 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[24]), 
          .D0(frac_add_Norm1[24]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[25]), 
          .D1(frac_add_Norm1[25]), .CIN(n61513), .S0(frac_Norm2[21]), 
          .S1(frac_Norm2[22]));
    defparam add_72_23.INIT0 = 16'hf690;
    defparam add_72_23.INIT1 = 16'hf690;
    defparam add_72_23.INJECT1_0 = "NO";
    defparam add_72_23.INJECT1_1 = "NO";
    LUT4 i12_2_lut (.A(frac[9]), .B(frac[14]), .Z(n37)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12_2_lut.init = 16'h8888;
    LUT4 i14_4_lut_adj_800 (.A(frac[19]), .B(frac[25]), .C(frac[24]), 
         .D(frac[6]), .Z(n39_adj_437)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i14_4_lut_adj_800.init = 16'h8000;
    LUT4 i9_2_lut_adj_801 (.A(frac[15]), .B(frac[20]), .Z(n34_adj_438)) /* synthesis lut_function=(A (B)) */ ;
    defparam i9_2_lut_adj_801.init = 16'h8888;
    CCU2D add_72_21 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[22]), 
          .D0(frac_add_Norm1[22]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[23]), 
          .D1(frac_add_Norm1[23]), .CIN(n61512), .COUT(n61513), .S0(frac_Norm2[19]), 
          .S1(frac_Norm2[20]));
    defparam add_72_21.INIT0 = 16'hf690;
    defparam add_72_21.INIT1 = 16'hf690;
    defparam add_72_21.INJECT1_0 = "NO";
    defparam add_72_21.INJECT1_1 = "NO";
    LUT4 i16_4_lut_adj_802 (.A(frac[13]), .B(frac[18]), .C(frac[22]), 
         .D(frac[23]), .Z(n41)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut_adj_802.init = 16'h8000;
    LUT4 i20_4_lut (.A(n39_adj_437), .B(frac[17]), .C(n30), .D(n70707), 
         .Z(n45)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_803 (.A(expB_FF), .B(expA_FF), .C(n66192), .D(n66206), 
         .Z(n4_adj_439)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_803.init = 16'heca0;
    LUT4 i19_4_lut_adj_804 (.A(n37), .B(frac[10]), .C(frac[7]), .D(frac[8]), 
         .Z(n44_adj_440)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19_4_lut_adj_804.init = 16'h8000;
    LUT4 i23_4_lut (.A(n45), .B(n41), .C(n33), .D(n34_adj_438), .Z(n48)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23_4_lut.init = 16'h8000;
    LUT4 i18_4_lut_adj_805 (.A(n70714), .B(frac[16]), .C(frac[12]), .D(frac[21]), 
         .Z(n43)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18_4_lut_adj_805.init = 16'h8000;
    LUT4 i63_4_lut (.A(frac[27]), .B(n43), .C(n48), .D(n44_adj_440), 
         .Z(n574)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i63_4_lut.init = 16'heaaa;
    CCU2D add_72_19 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[20]), 
          .D0(frac_add_Norm1[20]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[21]), 
          .D1(frac_add_Norm1[21]), .CIN(n61511), .COUT(n61512), .S0(frac_Norm2[17]), 
          .S1(frac_Norm2[18]));
    defparam add_72_19.INIT0 = 16'hf690;
    defparam add_72_19.INIT1 = 16'hf690;
    defparam add_72_19.INJECT1_0 = "NO";
    defparam add_72_19.INJECT1_1 = "NO";
    CCU2D add_72_17 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[18]), 
          .D0(frac_add_Norm1[18]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[19]), 
          .D1(frac_add_Norm1[19]), .CIN(n61510), .COUT(n61511), .S0(frac_Norm2[15]), 
          .S1(frac_Norm2[16]));
    defparam add_72_17.INIT0 = 16'hf690;
    defparam add_72_17.INIT1 = 16'hf690;
    defparam add_72_17.INJECT1_0 = "NO";
    defparam add_72_17.INJECT1_1 = "NO";
    CCU2D add_72_15 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[16]), 
          .D0(frac_add_Norm1[16]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[17]), 
          .D1(frac_add_Norm1[17]), .CIN(n61509), .COUT(n61510), .S0(frac_Norm2[13]), 
          .S1(frac_Norm2[14]));
    defparam add_72_15.INIT0 = 16'hf690;
    defparam add_72_15.INIT1 = 16'hf690;
    defparam add_72_15.INJECT1_0 = "NO";
    defparam add_72_15.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(expB_FF), .B(n4_adj_439), .C(n70805), .D(expA_FF), 
         .Z(n66234)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;
    defparam i2_4_lut.init = 16'hcecc;
    CCU2D add_72_13 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[14]), 
          .D0(frac_add_Norm1[14]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[15]), 
          .D1(frac_add_Norm1[15]), .CIN(n61508), .COUT(n61509), .S0(frac_Norm2[11]), 
          .S1(frac_Norm2[12]));
    defparam add_72_13.INIT0 = 16'hf690;
    defparam add_72_13.INIT1 = 16'hf690;
    defparam add_72_13.INJECT1_0 = "NO";
    defparam add_72_13.INJECT1_1 = "NO";
    CCU2D add_72_11 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[12]), 
          .D0(frac_add_Norm1[12]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[13]), 
          .D1(frac_add_Norm1[13]), .CIN(n61507), .COUT(n61508), .S0(frac_Norm2[9]), 
          .S1(frac_Norm2[10]));
    defparam add_72_11.INIT0 = 16'hf690;
    defparam add_72_11.INIT1 = 16'hf690;
    defparam add_72_11.INJECT1_0 = "NO";
    defparam add_72_11.INJECT1_1 = "NO";
    LUT4 mux_216_i6_3_lut (.A(n70703), .B(frac[6]), .C(frac[27]), .Z(frac_add_Norm1[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i6_3_lut.init = 16'hcaca;
    LUT4 mux_216_i5_3_lut (.A(n70706), .B(n70703), .C(frac[27]), .Z(frac_add_Norm1[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i5_3_lut.init = 16'hcaca;
    LUT4 mux_216_i8_3_lut (.A(frac[7]), .B(frac[8]), .C(frac[27]), .Z(frac_add_Norm1[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i8_3_lut.init = 16'hcaca;
    LUT4 mux_216_i7_3_lut (.A(frac[6]), .B(frac[7]), .C(frac[27]), .Z(frac_add_Norm1[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i7_3_lut.init = 16'hcaca;
    LUT4 mux_216_i10_3_lut (.A(frac[9]), .B(frac[10]), .C(frac[27]), .Z(frac_add_Norm1[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i10_3_lut.init = 16'hcaca;
    LUT4 mux_216_i9_3_lut (.A(frac[8]), .B(frac[9]), .C(frac[27]), .Z(frac_add_Norm1[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i9_3_lut.init = 16'hcaca;
    LUT4 mux_216_i12_3_lut (.A(frac[11]), .B(frac[12]), .C(frac[27]), 
         .Z(frac_add_Norm1[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i12_3_lut.init = 16'hcaca;
    CCU2D add_72_9 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[10]), 
          .D0(frac_add_Norm1[10]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[11]), 
          .D1(frac_add_Norm1[11]), .CIN(n61506), .COUT(n61507), .S0(frac_Norm2[7]), 
          .S1(frac_Norm2[8]));
    defparam add_72_9.INIT0 = 16'hf690;
    defparam add_72_9.INIT1 = 16'hf690;
    defparam add_72_9.INJECT1_0 = "NO";
    defparam add_72_9.INJECT1_1 = "NO";
    LUT4 mux_216_i11_3_lut (.A(frac[10]), .B(frac[11]), .C(frac[27]), 
         .Z(frac_add_Norm1[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i11_3_lut.init = 16'hcaca;
    CCU2D add_72_7 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[8]), 
          .D0(frac_add_Norm1[8]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[9]), 
          .D1(frac_add_Norm1[9]), .CIN(n61505), .COUT(n61506), .S0(frac_Norm2[5]), 
          .S1(frac_Norm2[6]));
    defparam add_72_7.INIT0 = 16'hf690;
    defparam add_72_7.INIT1 = 16'hf690;
    defparam add_72_7.INJECT1_0 = "NO";
    defparam add_72_7.INJECT1_1 = "NO";
    LUT4 mux_216_i14_3_lut (.A(frac[13]), .B(frac[14]), .C(frac[27]), 
         .Z(frac_add_Norm1[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i14_3_lut.init = 16'hcaca;
    CCU2D add_72_5 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[6]), 
          .D0(frac_add_Norm1[6]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[7]), 
          .D1(frac_add_Norm1[7]), .CIN(n61504), .COUT(n61505), .S0(frac_Norm2[3]), 
          .S1(frac_Norm2[4]));
    defparam add_72_5.INIT0 = 16'hf690;
    defparam add_72_5.INIT1 = 16'hf690;
    defparam add_72_5.INJECT1_0 = "NO";
    defparam add_72_5.INJECT1_1 = "NO";
    LUT4 mux_216_i13_3_lut (.A(frac[12]), .B(frac[13]), .C(frac[27]), 
         .Z(frac_add_Norm1[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i13_3_lut.init = 16'hcaca;
    LUT4 mux_216_i16_3_lut (.A(frac[15]), .B(frac[16]), .C(frac[27]), 
         .Z(frac_add_Norm1[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i16_3_lut.init = 16'hcaca;
    CCU2D add_72_3 (.A0(n70865), .B0(A_int[31]), .C0(frac_sub_Norm1[4]), 
          .D0(frac_add_Norm1[4]), .A1(n70865), .B1(A_int[31]), .C1(frac_sub_Norm1[5]), 
          .D1(frac_add_Norm1[5]), .CIN(n61503), .COUT(n61504), .S0(frac_Norm2[1]), 
          .S1(frac_Norm2[2]));
    defparam add_72_3.INIT0 = 16'hf690;
    defparam add_72_3.INIT1 = 16'hf690;
    defparam add_72_3.INJECT1_0 = "NO";
    defparam add_72_3.INJECT1_1 = "NO";
    LUT4 mux_216_i15_3_lut (.A(frac[14]), .B(frac[15]), .C(frac[27]), 
         .Z(frac_add_Norm1[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i15_3_lut.init = 16'hcaca;
    LUT4 mux_216_i18_3_lut (.A(frac[17]), .B(frac[18]), .C(frac[27]), 
         .Z(frac_add_Norm1[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i18_3_lut.init = 16'hcaca;
    CCU2D add_72_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(frac_Norm1[3]), .B1(n63665), .C1(n63661), .D1(frac_Norm1[2]), 
          .COUT(n61503), .S1(frac_Norm2[0]));
    defparam add_72_1.INIT0 = 16'hF000;
    defparam add_72_1.INIT1 = 16'h56a6;
    defparam add_72_1.INJECT1_0 = "NO";
    defparam add_72_1.INJECT1_1 = "NO";
    LUT4 mux_216_i17_3_lut (.A(frac[16]), .B(frac[17]), .C(frac[27]), 
         .Z(frac_add_Norm1[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i17_3_lut.init = 16'hcaca;
    LUT4 mux_216_i20_3_lut (.A(frac[19]), .B(frac[20]), .C(frac[27]), 
         .Z(frac_add_Norm1[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i20_3_lut.init = 16'hcaca;
    LUT4 mux_216_i19_3_lut (.A(frac[18]), .B(frac[19]), .C(frac[27]), 
         .Z(frac_add_Norm1[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i19_3_lut.init = 16'hcaca;
    LUT4 mux_216_i22_3_lut (.A(frac[21]), .B(frac[22]), .C(frac[27]), 
         .Z(frac_add_Norm1[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i22_3_lut.init = 16'hcaca;
    LUT4 mux_216_i21_3_lut (.A(frac[20]), .B(frac[21]), .C(frac[27]), 
         .Z(frac_add_Norm1[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i21_3_lut.init = 16'hcaca;
    LUT4 mux_216_i24_3_lut (.A(frac[23]), .B(frac[24]), .C(frac[27]), 
         .Z(frac_add_Norm1[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i24_3_lut.init = 16'hcaca;
    LUT4 mux_216_i23_3_lut (.A(frac[22]), .B(frac[23]), .C(frac[27]), 
         .Z(frac_add_Norm1[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i23_3_lut.init = 16'hcaca;
    LUT4 mux_216_i26_3_lut (.A(frac[25]), .B(frac[26]), .C(frac[27]), 
         .Z(frac_add_Norm1[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i26_3_lut.init = 16'hcaca;
    LUT4 mux_216_i25_3_lut (.A(frac[24]), .B(frac[25]), .C(frac[27]), 
         .Z(frac_add_Norm1[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_216_i25_3_lut.init = 16'hcaca;
    LUT4 mux_3773_i21_4_lut (.A(frac_Norm2[20]), .B(frac[23]), .C(n70739), 
         .D(n70613), .Z(n10673[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i21_4_lut.init = 16'hcac0;
    LUT4 i4_2_lut (.A(n8360[5]), .B(n8360[1]), .Z(n13_adj_441)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4_2_lut.init = 16'h8888;
    LUT4 i29915_2_lut_3_lut_4_lut (.A(B_int[31]), .B(add_enable), .C(leadZerosBin[1]), 
         .D(A_int[31]), .Z(n41510)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i29915_2_lut_3_lut_4_lut.init = 16'hf9f6;
    LUT4 i29911_2_lut_3_lut_4_lut (.A(B_int[31]), .B(add_enable), .C(n73795), 
         .D(A_int[31]), .Z(n41506)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i29911_2_lut_3_lut_4_lut.init = 16'hf9f6;
    LUT4 i29913_2_lut_3_lut_4_lut (.A(B_int[31]), .B(add_enable), .C(leadZerosBin[2]), 
         .D(A_int[31]), .Z(n41508)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i29913_2_lut_3_lut_4_lut.init = 16'hf9f6;
    LUT4 i6697_4_lut_3_lut_4_lut (.A(B_int[31]), .B(add_enable), .C(n17318), 
         .D(A_int[31]), .Z(sign)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i6697_4_lut_3_lut_4_lut.init = 16'h9f90;
    LUT4 i10006_1_lut_2_lut_3_lut (.A(B_int[31]), .B(add_enable), .C(A_int[31]), 
         .Z(isSUB)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam i10006_1_lut_2_lut_3_lut.init = 16'h6969;
    LUT4 i1_2_lut_rep_835_3_lut (.A(B_int[31]), .B(add_enable), .C(A_int[31]), 
         .Z(n70805)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_2_lut_rep_835_3_lut.init = 16'h9696;
    LUT4 i5097_2_lut_rep_895 (.A(B_int[31]), .B(add_enable), .Z(n70865)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5097_2_lut_rep_895.init = 16'h6666;
    LUT4 i1_4_lut_adj_806 (.A(n41778), .B(n70805), .C(\diffExp[4] ), .D(n7), 
         .Z(n21669)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_806.init = 16'hccc6;
    LUT4 i7_4_lut_adj_807 (.A(n13_adj_441), .B(n8360[7]), .C(n8360[0]), 
         .D(n41758), .Z(n16)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_807.init = 16'h8000;
    LUT4 i6_4_lut_adj_808 (.A(n8360[6]), .B(n8360[4]), .C(n8360[2]), .D(n8360[3]), 
         .Z(n15_adj_442)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut_adj_808.init = 16'h8000;
    LUT4 i1_4_lut_adj_809 (.A(n70777), .B(n70805), .C(n41588), .D(n7), 
         .Z(n21679)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_809.init = 16'hcc9c;
    LUT4 i1_4_lut_adj_810 (.A(n15_adj_443), .B(n70805), .C(n7), .D(n70743), 
         .Z(n21645)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_810.init = 16'hccc6;
    LUT4 i1_4_lut_adj_811 (.A(n7), .B(n70805), .C(n66914), .D(diffExp[2]), 
         .Z(n21651)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_811.init = 16'hcc9c;
    LUT4 i1_4_lut_adj_812 (.A(n7), .B(n70805), .C(n66904), .D(n70832), 
         .Z(n21643)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_812.init = 16'hcc9c;
    LUT4 i2_4_lut_adj_813 (.A(expB_FF), .B(n15_adj_442), .C(expA_FF), 
         .D(n16), .Z(n22565)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_813.init = 16'heca0;
    LUT4 i30174_2_lut_4_lut (.A(n53), .B(n70805), .C(n62965), .D(n41758), 
         .Z(n40687)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i30174_2_lut_4_lut.init = 16'hec00;
    LUT4 i1_4_lut_adj_814 (.A(expA_FF), .B(n70805), .C(expB_FF), .D(n22565), 
         .Z(n731)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_814.init = 16'hde5a;
    LUT4 mux_3773_i20_4_lut (.A(frac_Norm2[19]), .B(frac[22]), .C(n70739), 
         .D(n70613), .Z(n10673[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3773_i20_4_lut.init = 16'hcac0;
    LUT4 i12459_3_lut (.A(n73803), .B(n731), .C(n66234), .Z(n24122)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i12459_3_lut.init = 16'ha8a8;
    CCU2D add_3798_9 (.A0(n70805), .B0(A_int[29]), .C0(B_int[29]), .D0(diffExpAB[8]), 
          .A1(n70805), .B1(A_int[30]), .C1(B_int[30]), .D1(diffExpAB[8]), 
          .CIN(n61613), .S0(n8360[6]), .S1(n8360[7]));
    defparam add_3798_9.INIT0 = 16'ha599;
    defparam add_3798_9.INIT1 = 16'ha599;
    defparam add_3798_9.INJECT1_0 = "NO";
    defparam add_3798_9.INJECT1_1 = "NO";
    CCU2D add_3798_7 (.A0(n40002), .B0(A_int[27]), .C0(B_int[27]), .D0(diffExpAB[8]), 
          .A1(n70805), .B1(A_int[28]), .C1(B_int[28]), .D1(diffExpAB[8]), 
          .CIN(n61612), .COUT(n61613), .S0(n8360[4]), .S1(n8360[5]));
    defparam add_3798_7.INIT0 = 16'ha599;
    defparam add_3798_7.INIT1 = 16'ha599;
    defparam add_3798_7.INJECT1_0 = "NO";
    defparam add_3798_7.INJECT1_1 = "NO";
    CCU2D add_3798_5 (.A0(n41508), .B0(A_int[25]), .C0(B_int[25]), .D0(diffExpAB[8]), 
          .A1(n41506), .B1(A_int[26]), .C1(B_int[26]), .D1(diffExpAB[8]), 
          .CIN(n61611), .COUT(n61612), .S0(n8360[2]), .S1(n8360[3]));
    defparam add_3798_5.INIT0 = 16'ha599;
    defparam add_3798_5.INIT1 = 16'ha599;
    defparam add_3798_5.INJECT1_0 = "NO";
    defparam add_3798_5.INJECT1_1 = "NO";
    LUT4 i6853_2_lut_rep_653_3_lut_4_lut (.A(n70638), .B(n70726), .C(leadZerosBin[2]), 
         .D(n73795), .Z(n70623)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i6853_2_lut_rep_653_3_lut_4_lut.init = 16'hfffd;
    LUT4 mux_52_i9_3_lut (.A(A_int[5]), .B(B_int[5]), .C(n70737), .Z(n480[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i9_3_lut.init = 16'hacac;
    CCU2D add_3798_3 (.A0(efectExp[0]), .B0(leadZerosBin[0]), .C0(n574), 
          .D0(n70805), .A1(n41510), .B1(A_int[24]), .C1(B_int[24]), 
          .D1(diffExpAB[8]), .CIN(n61610), .COUT(n61611), .S0(n8360[0]), 
          .S1(n8360[1]));
    defparam add_3798_3.INIT0 = 16'h5a99;
    defparam add_3798_3.INIT1 = 16'ha599;
    defparam add_3798_3.INJECT1_0 = "NO";
    defparam add_3798_3.INJECT1_1 = "NO";
    CCU2D add_3798_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(A_int[31]), .B1(n70865), .C1(GND_net), .D1(GND_net), .COUT(n61610));
    defparam add_3798_1.INIT0 = 16'hF000;
    defparam add_3798_1.INIT1 = 16'h6666;
    defparam add_3798_1.INJECT1_0 = "NO";
    defparam add_3798_1.INJECT1_1 = "NO";
    LUT4 mux_51_i9_3_lut (.A(addSubAB[8]), .B(subBAExpEq[8]), .C(n70733), 
         .Z(n451[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i9_3_lut.init = 16'hcaca;
    LUT4 mux_52_i8_3_lut (.A(\A_int[4] ), .B(\B_int[4] ), .C(n70737), 
         .Z(n480[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i8_3_lut.init = 16'hacac;
    LUT4 mux_51_i8_3_lut (.A(addSubAB[7]), .B(subBAExpEq[7]), .C(n70733), 
         .Z(n451[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i8_3_lut.init = 16'hcaca;
    LUT4 mux_52_i11_3_lut (.A(\A_int[7] ), .B(\B_int[7] ), .C(n70737), 
         .Z(n480[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i11_3_lut.init = 16'hacac;
    LUT4 mux_51_i11_3_lut (.A(addSubAB[10]), .B(subBAExpEq[10]), .C(n70733), 
         .Z(n451[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i11_3_lut.init = 16'hcaca;
    LUT4 mux_52_i10_3_lut (.A(A_int[6]), .B(B_int[6]), .C(n70737), .Z(n480[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i10_3_lut.init = 16'hacac;
    LUT4 mux_51_i10_3_lut (.A(addSubAB[9]), .B(subBAExpEq[9]), .C(n70733), 
         .Z(n451[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_51_i10_3_lut.init = 16'hcaca;
    LUT4 mux_52_i13_3_lut (.A(\A_int[9] ), .B(\B_int[9] ), .C(n70737), 
         .Z(n480[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_52_i13_3_lut.init = 16'hacac;
    \fp_leading_zeros_and_shift(27,8,4)_U26  subtraction_norm (.n31(n31_adj_423), 
            .\leadZerosBin[2] (leadZerosBin[2]), .\leadZerosBin[1] (leadZerosBin[1]), 
            .\addSubAB[0] (addSubAB[0]), .n70638(n70638), .\efectExp[4] (efectExp[4]), 
            .\frac[21] (frac[21]), .n70703(n70703), .\frac[20] (frac[20]), 
            .n70706(n70706), .\frac[19] (frac[19]), .n70707(n70707), .\frac[11] (frac[11]), 
            .n73795(n73795), .n19138(n19138), .\frac[15] (frac[15]), .\frac[23] (frac[23]), 
            .\frac[7] (frac[7]), .\frac[14] (frac[14]), .\frac[22] (frac[22]), 
            .\frac[6] (frac[6]), .\addSubAB[1] (addSubAB[1]), .n70633(n70633), 
            .n70726(n70726), .\efectExp[0] (efectExp[0]), .\efectExp[1] (efectExp[1]), 
            .\leadZerosBin[0] (leadZerosBin[0]), .n19(n19), .\frac_sub_Norm1[4] (frac_sub_Norm1[4]), 
            .n70623(n70623), .n356(n330[2]), .\addSubAB[27] (addSubAB[27]), 
            .\subBAExpEq[27] (subBAExpEq[27]), .n70733(n70733), .\frac[27] (frac[27]), 
            .n21808(n21808), .\frac[10] (frac[10]), .\frac[16] (frac[16]), 
            .\frac[17] (frac[17]), .\frac[18] (frac[18]), .\frac[25] (frac[25]), 
            .\frac[26] (frac[26]), .\frac[24] (frac[24]), .n70641(n70641), 
            .n70643(n70643), .n39(n39), .n53(n53), .n70715(n70715), 
            .n70714(n70714), .\A_int[26] (A_int[26]), .\B_int[26] (B_int[26]), 
            .\diffExpAB[8] (diffExpAB[8]), .n70784(n70784), .\frac_sub_Norm1[3] (frac_sub_Norm1[3]), 
            .n70739(n70739), .\A_int[25] (A_int[25]), .\B_int[25] (B_int[25]), 
            .\efectExp[2] (efectExp[2]), .\A_int[24] (A_int[24]), .\B_int[24] (B_int[24]), 
            .\addSubAB[26] (addSubAB[26]), .\subBAExpEq[26] (subBAExpEq[26]), 
            .\frac[8] (frac[8]), .\frac[12] (frac[12]), .\frac[13] (frac[13]), 
            .n66182(n66182), .\frac_sub_Norm1[25] (frac_sub_Norm1[25]), 
            .n67677(n67677), .n66192(n66192), .n13(n13), .n14(n14_adj_436), 
            .\frac[9] (frac[9]), .\A_int[23] (A_int[23]), .\B_int[23] (B_int[23]), 
            .n70637(n70637), .\addSubAB[2] (addSubAB[2]), .n70636(n70636), 
            .n23602(n23602), .n66558(n66558), .n19142(n19142), .n19140(n19140), 
            .\frac_add_Norm1[2] (frac_add_Norm1[2]), .n476(n451[3]), .n505(n480[3]), 
            .n24(n24), .n475(n451[4]), .n504(n480[4]), .n25(n25), .n33(n33), 
            .n474(n451[5]), .n503(n480[5]), .n30(n30), .\A_int[27] (A_int[27]), 
            .\B_int[27] (B_int[27]), .\A_int[28] (A_int[28]), .\B_int[28] (B_int[28]), 
            .\efectExp[5] (efectExp[5]), .n266(n243[5]), .n291(n272[9]), 
            .n290(n272[10]), .n289(n272[11]), .n261(n243[10]), .n260(n243[11]), 
            .n259(n243[12]), .n258(n243[13]), .\A_int[29] (A_int[29]), 
            .\B_int[29] (B_int[29]), .\efectExp[6] (efectExp[6]), .\A_int[30] (A_int[30]), 
            .\B_int[30] (B_int[30]), .\efectExp[7] (efectExp[7]), .n454(n451[25]), 
            .n483(n480[25]), .n456(n451[23]), .n485(n480[23]), .n455(n451[24]), 
            .n484(n480[24]), .n458(n451[21]), .n487(n480[21]), .n457(n451[22]), 
            .n486(n480[22]), .n460(n451[19]), .n489(n480[19]), .n459(n451[20]), 
            .n488(n480[20]), .n462(n451[17]), .n491(n480[17]), .n461(n451[18]), 
            .n490(n480[18]), .n464(n451[15]), .n493(n480[15]), .n463(n451[16]), 
            .n492(n480[16]), .n466(n451[13]), .n495(n480[13]), .n465(n451[14]), 
            .n494(n480[14]), .n468(n451[11]), .n497(n480[11]), .n467(n451[12]), 
            .n496(n480[12]), .n470(n451[9]), .n499(n480[9]), .n469(n451[10]), 
            .n498(n480[10]), .n472(n451[7]), .n501(n480[7]), .n471(n451[8]), 
            .n500(n480[8]), .n62965(n62965), .\frac_sub_Norm1[5] (frac_sub_Norm1[5]), 
            .n4(n4), .\frac_sub_Norm1[7] (frac_sub_Norm1[7]), .\frac_sub_Norm1[6] (frac_sub_Norm1[6]), 
            .n265(n243[6]), .\frac_sub_Norm1[9] (frac_sub_Norm1[9]), .\frac_sub_Norm1[8] (frac_sub_Norm1[8]), 
            .\frac_sub_Norm1[11] (frac_sub_Norm1[11]), .\frac_sub_Norm1[10] (frac_sub_Norm1[10]), 
            .\frac_sub_Norm1[13] (frac_sub_Norm1[13]), .\frac_sub_Norm1[12] (frac_sub_Norm1[12]), 
            .n263(n243[8]), .\frac_sub_Norm1[15] (frac_sub_Norm1[15]), .\frac_sub_Norm1[14] (frac_sub_Norm1[14]), 
            .\frac_sub_Norm1[17] (frac_sub_Norm1[17]), .\frac_sub_Norm1[16] (frac_sub_Norm1[16]), 
            .\frac_sub_Norm1[19] (frac_sub_Norm1[19]), .\frac_sub_Norm1[18] (frac_sub_Norm1[18]), 
            .\frac_sub_Norm1[21] (frac_sub_Norm1[21]), .\frac_sub_Norm1[20] (frac_sub_Norm1[20]), 
            .\frac_sub_Norm1[23] (frac_sub_Norm1[23]), .\frac_sub_Norm1[22] (frac_sub_Norm1[22]), 
            .\frac_sub_Norm1[24] (frac_sub_Norm1[24]), .n66653(n66653), 
            .n17(n17), .\addSubAB[6] (addSubAB[6]), .\subBAExpEq[6] (subBAExpEq[6]), 
            .\B_int[3] (\B_int[3] ), .\A_int[3] (\A_int[3] ), .n70737(n70737), 
            .\frac_sub_Norm1[2] (frac_sub_Norm1[2]));
    \right_shifter(27,8,4)_U27  alignment (.diffExpAB({diffExpAB[8], diffExpAB_c[7:0]}), 
            .diffExpBA({diffExpBA}), .\diffExp[4] (\diffExp[4] ), .n70777(n70777), 
            .n70835(n70835), .\B_int[19] (B_int[19]), .\A_int[19] (A_int[19]), 
            .n70834(n70834), .\B_int[15] (B_int[15]), .\A_int[15] (A_int[15]), 
            .n70833(n70833), .n70832(n70832), .\B_int[1] (B_int[1]), .\A_int[1] (A_int[1]), 
            .\diffExp[2] (diffExp[2]), .\efectFracB[21] (\efectFracB[21] ), 
            .\efectFracB[20] (\efectFracB[20] ), .n70743(n70743), .\efectFracB[19] (\efectFracB[19] ), 
            .\efectFracB[15] (\efectFracB[15] ), .\efectFracB[16] (\efectFracB[16] ), 
            .n19214(n19214), .n15(n15_adj_443), .n28(n28), .n66904(n66904), 
            .n70771(n70771), .n9(n9), .\efectFracB[14] (\efectFracB[14] ), 
            .\efectFracB[7] (\efectFracB[7] ), .\efectFracB[5] (\efectFracB[5] ), 
            .\efectFracB[12] (\efectFracB[12] ), .n70820(n70820), .\efectFracB[13] (\efectFracB[13] ), 
            .n27(n27), .\fracAlign_int[0] (fracAlign_int[0]), .n70740(n70740), 
            .n7(n7), .\efectFracB_align[2] (efectFracB_align[2]), .\efectFracB_align[1] (efectFracB_align[1]), 
            .\B_int[0] (B_int[0]), .\A_int[0] (A_int[0]), .\fracAlign_int[4] (fracAlign_int[4]), 
            .\fracAlign_int[3] (fracAlign_int[3]), .n55(n55), .\fracAlign_int[6] (fracAlign_int[6]), 
            .\fracAlign_int[5] (fracAlign_int[5]), .\B_int[5] (B_int[5]), 
            .\A_int[5] (A_int[5]), .\fracAlign_int[8] (fracAlign_int[8]), 
            .\fracAlign_int[7] (fracAlign_int[7]), .\B_int[6] (B_int[6]), 
            .\A_int[6] (A_int[6]), .\fracAlign_int[10] (fracAlign_int[10]), 
            .\fracAlign_int[9] (fracAlign_int[9]), .\B_int[8] (B_int[8]), 
            .\A_int[8] (A_int[8]), .\fracAlign_int[12] (fracAlign_int[12]), 
            .n41778(n41778), .\fracAlign_int[14] (fracAlign_int[14]), .\fracAlign_int[13] (fracAlign_int[13]), 
            .\fracAlign_int[16] (fracAlign_int[16]), .\fracAlign_int[15] (fracAlign_int[15]), 
            .\fracAlign_int[18] (fracAlign_int[18]), .\fracAlign_int[17] (fracAlign_int[17]), 
            .\fracAlign_int[20] (fracAlign_int[20]), .n41588(n41588), .\fracAlign_int[22] (fracAlign_int[22]), 
            .\fracAlign_int[21] (fracAlign_int[21]), .n66914(n66914), .n66178(n66178), 
            .\B_int[22] (B_int[22]), .\A_int[22] (A_int[22]), .\B_int[14] (B_int[14]), 
            .\A_int[14] (A_int[14]), .\B_int[21] (B_int[21]), .\A_int[21] (A_int[21]), 
            .\B_int[20] (B_int[20]), .\A_int[20] (A_int[20]));
    
endmodule
//
// Verilog Description of module \fp_leading_zeros_and_shift(27,8,4)_U26 
//

module \fp_leading_zeros_and_shift(27,8,4)_U26  (n31, \leadZerosBin[2] , 
            \leadZerosBin[1] , \addSubAB[0] , n70638, \efectExp[4] , 
            \frac[21] , n70703, \frac[20] , n70706, \frac[19] , n70707, 
            \frac[11] , n73795, n19138, \frac[15] , \frac[23] , \frac[7] , 
            \frac[14] , \frac[22] , \frac[6] , \addSubAB[1] , n70633, 
            n70726, \efectExp[0] , \efectExp[1] , \leadZerosBin[0] , 
            n19, \frac_sub_Norm1[4] , n70623, n356, \addSubAB[27] , 
            \subBAExpEq[27] , n70733, \frac[27] , n21808, \frac[10] , 
            \frac[16] , \frac[17] , \frac[18] , \frac[25] , \frac[26] , 
            \frac[24] , n70641, n70643, n39, n53, n70715, n70714, 
            \A_int[26] , \B_int[26] , \diffExpAB[8] , n70784, \frac_sub_Norm1[3] , 
            n70739, \A_int[25] , \B_int[25] , \efectExp[2] , \A_int[24] , 
            \B_int[24] , \addSubAB[26] , \subBAExpEq[26] , \frac[8] , 
            \frac[12] , \frac[13] , n66182, \frac_sub_Norm1[25] , n67677, 
            n66192, n13, n14, \frac[9] , \A_int[23] , \B_int[23] , 
            n70637, \addSubAB[2] , n70636, n23602, n66558, n19142, 
            n19140, \frac_add_Norm1[2] , n476, n505, n24, n475, 
            n504, n25, n33, n474, n503, n30, \A_int[27] , \B_int[27] , 
            \A_int[28] , \B_int[28] , \efectExp[5] , n266, n291, n290, 
            n289, n261, n260, n259, n258, \A_int[29] , \B_int[29] , 
            \efectExp[6] , \A_int[30] , \B_int[30] , \efectExp[7] , 
            n454, n483, n456, n485, n455, n484, n458, n487, 
            n457, n486, n460, n489, n459, n488, n462, n491, 
            n461, n490, n464, n493, n463, n492, n466, n495, 
            n465, n494, n468, n497, n467, n496, n470, n499, 
            n469, n498, n472, n501, n471, n500, n62965, \frac_sub_Norm1[5] , 
            n4, \frac_sub_Norm1[7] , \frac_sub_Norm1[6] , n265, \frac_sub_Norm1[9] , 
            \frac_sub_Norm1[8] , \frac_sub_Norm1[11] , \frac_sub_Norm1[10] , 
            \frac_sub_Norm1[13] , \frac_sub_Norm1[12] , n263, \frac_sub_Norm1[15] , 
            \frac_sub_Norm1[14] , \frac_sub_Norm1[17] , \frac_sub_Norm1[16] , 
            \frac_sub_Norm1[19] , \frac_sub_Norm1[18] , \frac_sub_Norm1[21] , 
            \frac_sub_Norm1[20] , \frac_sub_Norm1[23] , \frac_sub_Norm1[22] , 
            \frac_sub_Norm1[24] , n66653, n17, \addSubAB[6] , \subBAExpEq[6] , 
            \B_int[3] , \A_int[3] , n70737, \frac_sub_Norm1[2] );
    output n31;
    input \leadZerosBin[2] ;
    output \leadZerosBin[1] ;
    input \addSubAB[0] ;
    input n70638;
    output \efectExp[4] ;
    output \frac[21] ;
    output n70703;
    output \frac[20] ;
    output n70706;
    output \frac[19] ;
    output n70707;
    output \frac[11] ;
    input n73795;
    output n19138;
    output \frac[15] ;
    output \frac[23] ;
    output \frac[7] ;
    output \frac[14] ;
    output \frac[22] ;
    output \frac[6] ;
    input \addSubAB[1] ;
    input n70633;
    input n70726;
    output \efectExp[0] ;
    output \efectExp[1] ;
    output \leadZerosBin[0] ;
    output n19;
    output \frac_sub_Norm1[4] ;
    input n70623;
    output n356;
    input \addSubAB[27] ;
    input \subBAExpEq[27] ;
    input n70733;
    output \frac[27] ;
    output n21808;
    output \frac[10] ;
    output \frac[16] ;
    output \frac[17] ;
    output \frac[18] ;
    output \frac[25] ;
    output \frac[26] ;
    output \frac[24] ;
    output n70641;
    output n70643;
    output n39;
    output n53;
    output n70715;
    output n70714;
    input \A_int[26] ;
    input \B_int[26] ;
    input \diffExpAB[8] ;
    output n70784;
    output \frac_sub_Norm1[3] ;
    output n70739;
    input \A_int[25] ;
    input \B_int[25] ;
    output \efectExp[2] ;
    input \A_int[24] ;
    input \B_int[24] ;
    input \addSubAB[26] ;
    input \subBAExpEq[26] ;
    output \frac[8] ;
    output \frac[12] ;
    output \frac[13] ;
    output n66182;
    output \frac_sub_Norm1[25] ;
    input n67677;
    input n66192;
    input n13;
    input n14;
    output \frac[9] ;
    input \A_int[23] ;
    input \B_int[23] ;
    input n70637;
    input \addSubAB[2] ;
    input n70636;
    input n23602;
    output n66558;
    output n19142;
    output n19140;
    output \frac_add_Norm1[2] ;
    input n476;
    input n505;
    output n24;
    input n475;
    input n504;
    output n25;
    output n33;
    input n474;
    input n503;
    output n30;
    input \A_int[27] ;
    input \B_int[27] ;
    input \A_int[28] ;
    input \B_int[28] ;
    output \efectExp[5] ;
    input n266;
    input n291;
    input n290;
    input n289;
    input n261;
    input n260;
    input n259;
    input n258;
    input \A_int[29] ;
    input \B_int[29] ;
    output \efectExp[6] ;
    input \A_int[30] ;
    input \B_int[30] ;
    output \efectExp[7] ;
    input n454;
    input n483;
    input n456;
    input n485;
    input n455;
    input n484;
    input n458;
    input n487;
    input n457;
    input n486;
    input n460;
    input n489;
    input n459;
    input n488;
    input n462;
    input n491;
    input n461;
    input n490;
    input n464;
    input n493;
    input n463;
    input n492;
    input n466;
    input n495;
    input n465;
    input n494;
    input n468;
    input n497;
    input n467;
    input n496;
    input n470;
    input n499;
    input n469;
    input n498;
    input n472;
    input n501;
    input n471;
    input n500;
    output n62965;
    output \frac_sub_Norm1[5] ;
    input n4;
    output \frac_sub_Norm1[7] ;
    output \frac_sub_Norm1[6] ;
    input n265;
    output \frac_sub_Norm1[9] ;
    output \frac_sub_Norm1[8] ;
    output \frac_sub_Norm1[11] ;
    output \frac_sub_Norm1[10] ;
    output \frac_sub_Norm1[13] ;
    output \frac_sub_Norm1[12] ;
    input n263;
    output \frac_sub_Norm1[15] ;
    output \frac_sub_Norm1[14] ;
    output \frac_sub_Norm1[17] ;
    output \frac_sub_Norm1[16] ;
    output \frac_sub_Norm1[19] ;
    output \frac_sub_Norm1[18] ;
    output \frac_sub_Norm1[21] ;
    output \frac_sub_Norm1[20] ;
    output \frac_sub_Norm1[23] ;
    output \frac_sub_Norm1[22] ;
    output \frac_sub_Norm1[24] ;
    output n66653;
    output n17;
    input \addSubAB[6] ;
    input \subBAExpEq[6] ;
    input \B_int[3] ;
    input \A_int[3] ;
    input n70737;
    output \frac_sub_Norm1[2] ;
    
    
    wire n24_c, n20, n18, n112, n114, n19_c, n70672, n70668, 
        n136, n70662, n23, n21, n138, n70671, n27, n121, n70632;
    wire [27:0]n330;
    
    wire n6, n8;
    wire [27:0]n243;
    wire [27:0]n272;
    
    wire n70616, n67113, n70630;
    wire [27:0]n301;
    
    wire n4_c, n19114, n70621, n70622, n67676, n5, n70646, n62779, 
        n66650, n22464, n9, n17_c, n10, n66680, n22, n22225, 
        n70663, n105, n70656, n66592, n35, n70650, n114_adj_412, 
        n22165, n49, n23588, n4_adj_413, n70130, n70629, n70127, 
        n70869, n70870, n70129, n70045, n70044, n66751, n66736, 
        n70043, n12, n70031, n70032, n70030, n70029, n70628, n70719, 
        n17316, n63537, n67170, n10_adj_415, n19122, n70685, n20408, 
        n19134, n20404, n19132, n19130, n70674;
    
    LUT4 i1_4_lut (.A(n24_c), .B(n20), .C(n18), .D(n112), .Z(n114)) /* synthesis lut_function=((B ((D)+!C))+!A) */ ;
    defparam i1_4_lut.init = 16'hdd5d;
    LUT4 i1_4_lut_adj_737 (.A(n19_c), .B(n70672), .C(n70668), .D(n114), 
         .Z(n136)) /* synthesis lut_function=(A ((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_737.init = 16'ha222;
    LUT4 i1_4_lut_adj_738 (.A(n70662), .B(n23), .C(n21), .D(n136), .Z(n138)) /* synthesis lut_function=((B ((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_738.init = 16'hdd5d;
    LUT4 i1_4_lut_adj_739 (.A(n31), .B(n70671), .C(n27), .D(n138), .Z(n121)) /* synthesis lut_function=(A ((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_739.init = 16'ha222;
    LUT4 i29150_3_lut_4_lut (.A(n70632), .B(\leadZerosBin[2] ), .C(\leadZerosBin[1] ), 
         .D(\addSubAB[0] ), .Z(n330[0])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i29150_3_lut_4_lut.init = 16'h0100;
    LUT4 LessThan_87_i8_3_lut_3_lut (.A(n70638), .B(\efectExp[4] ), .C(n6), 
         .Z(n8)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;
    defparam LessThan_87_i8_3_lut_3_lut.init = 16'he8e8;
    LUT4 mux_32_i22_3_lut (.A(\frac[21] ), .B(n70703), .C(n70638), .Z(n243[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_32_i22_3_lut.init = 16'hacac;
    LUT4 mux_32_i21_3_lut (.A(\frac[20] ), .B(n70706), .C(n70638), .Z(n243[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_32_i21_3_lut.init = 16'hacac;
    LUT4 mux_32_i20_3_lut (.A(\frac[19] ), .B(n70707), .C(n70638), .Z(n243[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_32_i20_3_lut.init = 16'hacac;
    LUT4 i7838_3_lut (.A(\frac[11] ), .B(n70707), .C(n73795), .Z(n19138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7838_3_lut.init = 16'hcaca;
    LUT4 mux_30_i24_4_lut (.A(\frac[15] ), .B(n272[19]), .C(\leadZerosBin[2] ), 
         .D(n70638), .Z(n272[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_30_i24_4_lut.init = 16'hcac0;
    LUT4 mux_32_i24_3_lut (.A(\frac[23] ), .B(\frac[7] ), .C(n70638), 
         .Z(n243[23])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_32_i24_3_lut.init = 16'hacac;
    LUT4 mux_30_i23_4_lut (.A(\frac[14] ), .B(n272[18]), .C(\leadZerosBin[2] ), 
         .D(n70638), .Z(n272[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_30_i23_4_lut.init = 16'hcac0;
    LUT4 mux_32_i23_3_lut (.A(\frac[22] ), .B(\frac[6] ), .C(n70638), 
         .Z(n243[22])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_32_i23_3_lut.init = 16'hacac;
    LUT4 i2_2_lut_rep_646_4_lut (.A(\addSubAB[1] ), .B(n70633), .C(n70726), 
         .D(\leadZerosBin[1] ), .Z(n70616)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_2_lut_rep_646_4_lut.init = 16'h0002;
    LUT4 mux_26_i5_3_lut_4_lut (.A(n67113), .B(n70630), .C(\leadZerosBin[1] ), 
         .D(n301[4]), .Z(n330[4])) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_26_i5_3_lut_4_lut.init = 16'h4f40;
    LUT4 LessThan_87_i4_4_lut (.A(\efectExp[0] ), .B(\efectExp[1] ), .C(\leadZerosBin[1] ), 
         .D(\leadZerosBin[0] ), .Z(n4_c)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;
    defparam LessThan_87_i4_4_lut.init = 16'h0c8e;
    LUT4 i1_3_lut_4_lut (.A(\leadZerosBin[2] ), .B(n70616), .C(n330[0]), 
         .D(\leadZerosBin[0] ), .Z(n19)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i55097_2_lut (.A(\leadZerosBin[2] ), .B(n73795), .Z(n67113)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i55097_2_lut.init = 16'heeee;
    LUT4 mux_21_i5_3_lut_4_lut (.A(n19114), .B(\leadZerosBin[2] ), .C(\leadZerosBin[0] ), 
         .D(n330[4]), .Z(\frac_sub_Norm1[4] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_21_i5_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_26_i3_4_lut (.A(n70621), .B(\addSubAB[0] ), .C(\leadZerosBin[1] ), 
         .D(n70623), .Z(n356)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_26_i3_4_lut.init = 16'h0aca;
    LUT4 i7814_4_lut (.A(n70707), .B(n70622), .C(\leadZerosBin[1] ), .D(n70633), 
         .Z(n19114)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam i7814_4_lut.init = 16'hc0ca;
    LUT4 i29458_4_lut (.A(\addSubAB[27] ), .B(n67676), .C(\subBAExpEq[27] ), 
         .D(n70733), .Z(\frac[27] )) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29458_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_740 (.A(n5), .B(n70646), .C(n62779), .D(n66650), 
         .Z(n21808)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_740.init = 16'h3b33;
    LUT4 i1_2_lut (.A(\frac[10] ), .B(n31), .Z(n22464)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 equal_58_i9_2_lut (.A(\frac[19] ), .B(\frac[20] ), .Z(n9)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_58_i9_2_lut.init = 16'heeee;
    LUT4 equal_40_i17_2_lut (.A(\frac[16] ), .B(\frac[17] ), .Z(n17_c)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_40_i17_2_lut.init = 16'heeee;
    LUT4 equal_55_i10_2_lut (.A(\frac[18] ), .B(\frac[19] ), .Z(n10)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_55_i10_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_741 (.A(\frac[15] ), .B(n21), .Z(n23)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_741.init = 16'heeee;
    LUT4 i3_4_lut (.A(\frac[18] ), .B(n17_c), .C(n9), .D(n20), .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_742 (.A(n19_c), .B(n21), .Z(n5)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_742.init = 16'h8888;
    LUT4 i1_2_lut_adj_743 (.A(\frac[21] ), .B(n18), .Z(n20)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_743.init = 16'heeee;
    LUT4 i1_2_lut_adj_744 (.A(\frac[20] ), .B(n66680), .Z(n24_c)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_744.init = 16'heeee;
    LUT4 equal_76_i3_2_lut (.A(\frac[25] ), .B(\frac[26] ), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_76_i3_2_lut.init = 16'heeee;
    LUT4 i2_4_lut (.A(\frac[24] ), .B(\frac[23] ), .C(n22), .D(\frac[22] ), 
         .Z(n18)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_745 (.A(\frac[23] ), .B(\frac[24] ), .Z(n22225)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_745.init = 16'heeee;
    LUT4 i1_4_lut_adj_746 (.A(n22225), .B(n70663), .C(n18), .D(n22), 
         .Z(n105)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A (B))) */ ;
    defparam i1_4_lut_adj_746.init = 16'h33b3;
    LUT4 i1_4_lut_adj_747 (.A(n105), .B(n70656), .C(n5), .D(n66650), 
         .Z(n66592)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;
    defparam i1_4_lut_adj_747.init = 16'h8c0c;
    LUT4 i1_4_lut_adj_748 (.A(n66592), .B(n35), .C(n31), .D(n70650), 
         .Z(n114_adj_412)) /* synthesis lut_function=(A ((C)+!B)+!A !(B ((D)+!C))) */ ;
    defparam i1_4_lut_adj_748.init = 16'hb3f3;
    LUT4 i1_4_lut_adj_749 (.A(n114_adj_412), .B(n70641), .C(n70643), .D(n39), 
         .Z(n22165)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;
    defparam i1_4_lut_adj_749.init = 16'h8c0c;
    LUT4 i2_4_lut_adj_750 (.A(n22165), .B(n53), .C(n70715), .D(n49), 
         .Z(\leadZerosBin[1] )) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i2_4_lut_adj_750.init = 16'hbbbf;
    LUT4 i1_4_lut_adj_751 (.A(n70715), .B(\addSubAB[0] ), .C(n70714), 
         .D(n23588), .Z(n4_adj_413)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+(D)))) */ ;
    defparam i1_4_lut_adj_751.init = 16'h0a3b;
    LUT4 i26_4_lut (.A(n70726), .B(n70130), .C(n70641), .D(n4_adj_413), 
         .Z(\leadZerosBin[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i26_4_lut.init = 16'hcfca;
    LUT4 LessThan_87_i7_2_lut_rep_659_4_lut (.A(\A_int[26] ), .B(\B_int[26] ), 
         .C(\diffExpAB[8] ), .D(n73795), .Z(n70629)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam LessThan_87_i7_2_lut_rep_659_4_lut.init = 16'h35ca;
    LUT4 mux_212_i4_3_lut_rep_814 (.A(\A_int[26] ), .B(\B_int[26] ), .C(\diffExpAB[8] ), 
         .Z(n70784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i4_3_lut_rep_814.init = 16'hcaca;
    LUT4 mux_21_i4_3_lut_4_lut (.A(n19114), .B(\leadZerosBin[2] ), .C(\leadZerosBin[0] ), 
         .D(n356), .Z(\frac_sub_Norm1[3] )) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;
    defparam mux_21_i4_3_lut_4_lut.init = 16'hf202;
    LUT4 frac_5__bdd_4_lut (.A(n70703), .B(\frac[6] ), .C(n70706), .D(\frac[7] ), 
         .Z(n70127)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam frac_5__bdd_4_lut.init = 16'hff23;
    PFUMX i56076 (.BLUT(n70869), .ALUT(n70870), .C0(n70739), .Z(\frac[6] ));
    PFUMX i55872 (.BLUT(n70129), .ALUT(n121), .C0(n22464), .Z(n70130));
    LUT4 i29396_2_lut_3_lut (.A(n70638), .B(n73795), .C(\frac[7] ), .Z(n272[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29396_2_lut_3_lut.init = 16'h2020;
    LUT4 mux_212_i3_3_lut (.A(\A_int[25] ), .B(\B_int[25] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i3_3_lut.init = 16'hcaca;
    LUT4 i29397_2_lut_3_lut (.A(n70638), .B(n73795), .C(\frac[6] ), .Z(n272[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29397_2_lut_3_lut.init = 16'h2020;
    LUT4 n70045_bdd_3_lut (.A(n70045), .B(n301[22]), .C(\leadZerosBin[1] ), 
         .Z(n330[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70045_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_212_i2_3_lut (.A(\A_int[24] ), .B(\B_int[24] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i2_3_lut.init = 16'hcaca;
    LUT4 n70044_bdd_3_lut (.A(n70044), .B(n272[20]), .C(\leadZerosBin[2] ), 
         .Z(n70045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70044_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_752 (.A(\frac[15] ), .B(\frac[14] ), .Z(n66751)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_752.init = 16'heeee;
    LUT4 i1_2_lut_adj_753 (.A(\frac[21] ), .B(\frac[20] ), .Z(n66736)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_753.init = 16'heeee;
    LUT4 i29459_4_lut (.A(\addSubAB[26] ), .B(n70739), .C(\subBAExpEq[26] ), 
         .D(n70733), .Z(\frac[26] )) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i29459_4_lut.init = 16'hfcee;
    PFUMX i55826 (.BLUT(n70043), .ALUT(n243[16]), .C0(n73795), .Z(n70044));
    LUT4 n255_bdd_3_lut_56431 (.A(n70638), .B(\frac[24] ), .C(\frac[8] ), 
         .Z(n70043)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n255_bdd_3_lut_56431.init = 16'hd8d8;
    LUT4 i5_4_lut (.A(\frac[26] ), .B(\frac[25] ), .C(\frac[22] ), .D(n66736), 
         .Z(n12)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(n66751), .B(n12), .C(\frac[12] ), .D(\frac[13] ), 
         .Z(n66182)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 n70031_bdd_3_lut (.A(n70031), .B(n301[23]), .C(\leadZerosBin[1] ), 
         .Z(n70032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70031_bdd_3_lut.init = 16'hcaca;
    LUT4 n70030_bdd_3_lut (.A(n70030), .B(n272[21]), .C(\leadZerosBin[2] ), 
         .Z(n70031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70030_bdd_3_lut.init = 16'hcaca;
    PFUMX i55820 (.BLUT(n70029), .ALUT(n243[17]), .C0(n73795), .Z(n70030));
    LUT4 n70032_bdd_3_lut (.A(n70032), .B(n330[24]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[25] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n70032_bdd_3_lut.init = 16'hcaca;
    LUT4 i55059_1_lut_4_lut (.A(n67677), .B(n66192), .C(n13), .D(n14), 
         .Z(n67676)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;
    defparam i55059_1_lut_4_lut.init = 16'h5554;
    LUT4 i55062_4_lut_rep_769 (.A(n67677), .B(n66192), .C(n13), .D(n14), 
         .Z(n70739)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;
    defparam i55062_4_lut_rep_769.init = 16'haaab;
    LUT4 n254_bdd_3_lut_56476 (.A(n70638), .B(\frac[25] ), .C(\frac[9] ), 
         .Z(n70029)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n254_bdd_3_lut_56476.init = 16'hd8d8;
    LUT4 mux_212_i1_3_lut (.A(\A_int[23] ), .B(\B_int[23] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i1_3_lut.init = 16'hcaca;
    LUT4 i29398_2_lut_3_lut (.A(n70638), .B(n73795), .C(n70703), .Z(n272[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29398_2_lut_3_lut.init = 16'h2020;
    LUT4 i29599_3_lut_rep_652_4_lut (.A(n70638), .B(n73795), .C(n70726), 
         .D(\addSubAB[1] ), .Z(n70622)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i29599_3_lut_rep_652_4_lut.init = 16'h0200;
    LUT4 i29399_2_lut_rep_658_3_lut (.A(n70638), .B(n73795), .C(n70706), 
         .Z(n70628)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i29399_2_lut_rep_658_3_lut.init = 16'h2020;
    LUT4 i2_2_lut_rep_651_3_lut_4_lut (.A(\leadZerosBin[2] ), .B(n73795), 
         .C(n70637), .D(\addSubAB[2] ), .Z(n70621)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_2_lut_rep_651_3_lut_4_lut.init = 16'h0100;
    LUT4 i29128_2_lut_rep_749_3_lut (.A(n70733), .B(n70739), .C(\addSubAB[0] ), 
         .Z(n70719)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29128_2_lut_rep_749_3_lut.init = 16'h1010;
    LUT4 i6692_2_lut_3_lut_4_lut (.A(n70733), .B(n70739), .C(\frac[27] ), 
         .D(\addSubAB[1] ), .Z(n17316)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i6692_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i29590_2_lut_rep_745_3_lut (.A(n70733), .B(n70739), .C(\addSubAB[1] ), 
         .Z(n70715)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29590_2_lut_rep_745_3_lut.init = 16'h1010;
    LUT4 i2_3_lut_4_lut (.A(n70733), .B(n70739), .C(n70638), .D(\addSubAB[1] ), 
         .Z(n63537)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i29588_2_lut_rep_744_3_lut (.A(n70733), .B(n70739), .C(\addSubAB[2] ), 
         .Z(n70714)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29588_2_lut_rep_744_3_lut.init = 16'h1010;
    LUT4 i55093_4_lut_4_lut (.A(n70636), .B(\efectExp[2] ), .C(\leadZerosBin[2] ), 
         .D(n70629), .Z(n67170)) /* synthesis lut_function=((B ((D)+!C)+!B (C+(D)))+!A) */ ;
    defparam i55093_4_lut_4_lut.init = 16'hff7d;
    LUT4 i29579_2_lut_rep_660_3_lut_4_lut (.A(n70733), .B(n70739), .C(\addSubAB[2] ), 
         .D(n70638), .Z(n70630)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i29579_2_lut_rep_660_3_lut_4_lut.init = 16'h1000;
    LUT4 i6851_2_lut_rep_662_3_lut_4_lut (.A(n70733), .B(n70739), .C(n73795), 
         .D(n70638), .Z(n70632)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i6851_2_lut_rep_662_3_lut_4_lut.init = 16'hfeff;
    LUT4 LessThan_87_i6_3_lut_3_lut (.A(n73795), .B(n70784), .C(\efectExp[2] ), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;
    defparam LessThan_87_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_4_lut_4_lut (.A(\addSubAB[0] ), .B(n70726), .C(n23602), .D(n17316), 
         .Z(n66558)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'hff32;
    LUT4 mux_32_i17_3_lut_4_lut (.A(\addSubAB[0] ), .B(n70726), .C(n70638), 
         .D(\frac[16] ), .Z(n243[16])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;
    defparam mux_32_i17_3_lut_4_lut.init = 16'hf202;
    LUT4 i2_4_lut_4_lut (.A(\addSubAB[0] ), .B(n70726), .C(n70641), .D(n23588), 
         .Z(n53)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i2_4_lut_4_lut.init = 16'hf3f2;
    LUT4 mux_32_i18_3_lut_4_lut (.A(\addSubAB[1] ), .B(n70726), .C(n70638), 
         .D(\frac[17] ), .Z(n243[17])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;
    defparam mux_32_i18_3_lut_4_lut.init = 16'hf202;
    LUT4 i7842_3_lut_4_lut (.A(\addSubAB[1] ), .B(n70726), .C(n73795), 
         .D(\frac[9] ), .Z(n19142)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i7842_3_lut_4_lut.init = 16'h2f20;
    LUT4 i7840_3_lut_4_lut (.A(\addSubAB[2] ), .B(n70726), .C(n73795), 
         .D(\frac[10] ), .Z(n19140)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i7840_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_216_i3_3_lut_4_lut (.A(\addSubAB[2] ), .B(n70726), .C(\frac[27] ), 
         .D(n70707), .Z(\frac_add_Norm1[2] )) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;
    defparam mux_216_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 mux_32_i19_3_lut_4_lut (.A(\addSubAB[2] ), .B(n70726), .C(n70638), 
         .D(\frac[18] ), .Z(n243[18])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;
    defparam mux_32_i19_3_lut_4_lut.init = 16'hf202;
    LUT4 i4_2_lut_4_lut (.A(n476), .B(n505), .C(n70739), .D(n70719), 
         .Z(n24)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i4_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_53_i4_3_lut_rep_737 (.A(n476), .B(n505), .C(n70739), .Z(n70707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i4_3_lut_rep_737.init = 16'hcaca;
    LUT4 i5_2_lut_4_lut (.A(n475), .B(n504), .C(n70739), .D(\frac[16] ), 
         .Z(n25)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i5_2_lut_4_lut.init = 16'hffca;
    LUT4 i8_2_lut_4_lut (.A(n475), .B(n504), .C(n70739), .D(\frac[11] ), 
         .Z(n33)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i8_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_53_i5_3_lut_rep_736 (.A(n475), .B(n504), .C(n70739), .Z(n70706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i5_3_lut_rep_736.init = 16'hcaca;
    LUT4 i5_2_lut_4_lut_adj_754 (.A(n474), .B(n503), .C(n70739), .D(\frac[26] ), 
         .Z(n30)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i5_2_lut_4_lut_adj_754.init = 16'hca00;
    LUT4 mux_53_i6_3_lut_rep_733 (.A(n474), .B(n503), .C(n70739), .Z(n70703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i6_3_lut_rep_733.init = 16'hcaca;
    LUT4 mux_212_i5_3_lut (.A(\A_int[27] ), .B(\B_int[27] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i5_3_lut.init = 16'hcaca;
    LUT4 i11902_2_lut (.A(\addSubAB[1] ), .B(\addSubAB[2] ), .Z(n23588)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11902_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_rep_701_4_lut (.A(n10), .B(n17_c), .C(n66182), .D(n22225), 
         .Z(n70671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_701_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_692_4_lut (.A(n10), .B(n17_c), .C(n24_c), .D(n66751), 
         .Z(n70662)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_692_4_lut.init = 16'hfffe;
    PFUMX LessThan_87_i10 (.BLUT(n4_c), .ALUT(n8), .C0(n67170), .Z(n10_adj_415));
    LUT4 mux_212_i6_3_lut (.A(\A_int[28] ), .B(\B_int[28] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i6_3_lut.init = 16'hcaca;
    PFUMX mux_28_i23 (.BLUT(n243[22]), .ALUT(n272[22]), .C0(n67113), .Z(n301[22]));
    PFUMX mux_28_i24 (.BLUT(n243[23]), .ALUT(n272[23]), .C0(n67113), .Z(n301[23]));
    PFUMX i7822 (.BLUT(n266), .ALUT(n63537), .C0(\leadZerosBin[2] ), .Z(n19122));
    PFUMX mux_28_i10 (.BLUT(n291), .ALUT(n272[5]), .C0(\leadZerosBin[2] ), 
          .Z(n301[9]));
    PFUMX mux_28_i11 (.BLUT(n290), .ALUT(n272[6]), .C0(\leadZerosBin[2] ), 
          .Z(n301[10]));
    PFUMX mux_28_i12 (.BLUT(n289), .ALUT(n272[7]), .C0(\leadZerosBin[2] ), 
          .Z(n301[11]));
    PFUMX mux_30_i19 (.BLUT(n243[18]), .ALUT(n261), .C0(n73795), .Z(n272[18]));
    PFUMX mux_30_i20 (.BLUT(n243[19]), .ALUT(n260), .C0(n73795), .Z(n272[19]));
    PFUMX mux_30_i21 (.BLUT(n243[20]), .ALUT(n259), .C0(n73795), .Z(n272[20]));
    PFUMX mux_30_i22 (.BLUT(n243[21]), .ALUT(n258), .C0(n73795), .Z(n272[21]));
    LUT4 mux_212_i7_3_lut (.A(\A_int[29] ), .B(\B_int[29] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i7_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_adj_755 (.A(n22), .B(n22225), .C(\frac[22] ), 
         .D(\frac[21] ), .Z(n66680)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_755.init = 16'hfffe;
    LUT4 mux_212_i8_3_lut (.A(\A_int[30] ), .B(\B_int[30] ), .C(\diffExpAB[8] ), 
         .Z(\efectExp[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_212_i8_3_lut.init = 16'hcaca;
    PFUMX mux_53_i26 (.BLUT(n454), .ALUT(n483), .C0(n70739), .Z(\frac[25] ));
    PFUMX mux_53_i24 (.BLUT(n456), .ALUT(n485), .C0(n70739), .Z(\frac[23] ));
    PFUMX mux_53_i25 (.BLUT(n455), .ALUT(n484), .C0(n70739), .Z(\frac[24] ));
    PFUMX mux_53_i22 (.BLUT(n458), .ALUT(n487), .C0(n70739), .Z(\frac[21] ));
    PFUMX mux_53_i23 (.BLUT(n457), .ALUT(n486), .C0(n70739), .Z(\frac[22] ));
    PFUMX mux_53_i20 (.BLUT(n460), .ALUT(n489), .C0(n70739), .Z(\frac[19] ));
    PFUMX mux_53_i21 (.BLUT(n459), .ALUT(n488), .C0(n70739), .Z(\frac[20] ));
    PFUMX mux_53_i18 (.BLUT(n462), .ALUT(n491), .C0(n70739), .Z(\frac[17] ));
    PFUMX mux_53_i19 (.BLUT(n461), .ALUT(n490), .C0(n70739), .Z(\frac[18] ));
    PFUMX mux_53_i16 (.BLUT(n464), .ALUT(n493), .C0(n70739), .Z(\frac[15] ));
    PFUMX mux_53_i17 (.BLUT(n463), .ALUT(n492), .C0(n70739), .Z(\frac[16] ));
    PFUMX mux_53_i14 (.BLUT(n466), .ALUT(n495), .C0(n70739), .Z(\frac[13] ));
    PFUMX mux_53_i15 (.BLUT(n465), .ALUT(n494), .C0(n70739), .Z(\frac[14] ));
    PFUMX mux_53_i12 (.BLUT(n468), .ALUT(n497), .C0(n70739), .Z(\frac[11] ));
    PFUMX mux_53_i13 (.BLUT(n467), .ALUT(n496), .C0(n70739), .Z(\frac[12] ));
    PFUMX mux_53_i10 (.BLUT(n470), .ALUT(n499), .C0(n70739), .Z(\frac[9] ));
    PFUMX mux_53_i11 (.BLUT(n469), .ALUT(n498), .C0(n70739), .Z(\frac[10] ));
    PFUMX mux_53_i8 (.BLUT(n472), .ALUT(n501), .C0(n70739), .Z(\frac[7] ));
    PFUMX mux_53_i9 (.BLUT(n471), .ALUT(n500), .C0(n70739), .Z(\frac[8] ));
    LUT4 i3_4_lut_adj_756 (.A(n10_adj_415), .B(\efectExp[7] ), .C(\efectExp[6] ), 
         .D(\efectExp[5] ), .Z(n62965)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_756.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n66736), .B(n10), .C(n18), .D(\frac[17] ), 
         .Z(n19_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_rep_702 (.A(n66736), .B(n10), .C(n18), .Z(n70672)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_702.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_757 (.A(n70685), .B(n22225), .C(n66182), .D(\frac[11] ), 
         .Z(n31)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_757.init = 16'hfffe;
    LUT4 i28000_2_lut_rep_680_4_lut (.A(n70685), .B(n22225), .C(n66182), 
         .D(n27), .Z(n70650)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i28000_2_lut_rep_680_4_lut.init = 16'hfe00;
    LUT4 mux_21_i6_3_lut (.A(n330[5]), .B(n330[4]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i6_3_lut.init = 16'hcaca;
    LUT4 mux_26_i6_4_lut (.A(n301[5]), .B(n67113), .C(\leadZerosBin[1] ), 
         .D(n4), .Z(n330[5])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_26_i6_4_lut.init = 16'h3a0a;
    LUT4 mux_28_i5_4_lut (.A(n70628), .B(\addSubAB[0] ), .C(\leadZerosBin[2] ), 
         .D(n70632), .Z(n301[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_28_i5_4_lut.init = 16'h0aca;
    LUT4 mux_26_i7_3_lut (.A(n301[6]), .B(n301[4]), .C(\leadZerosBin[1] ), 
         .Z(n330[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i7_3_lut.init = 16'hcaca;
    LUT4 mux_21_i8_3_lut (.A(n330[7]), .B(n330[6]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i8_3_lut.init = 16'hcaca;
    LUT4 mux_21_i7_3_lut (.A(n330[6]), .B(n330[5]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i7_3_lut.init = 16'hcaca;
    LUT4 i29387_2_lut (.A(n19122), .B(n73795), .Z(n301[5])) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i29387_2_lut.init = 16'h2222;
    LUT4 mux_26_i8_3_lut (.A(n301[7]), .B(n301[5]), .C(\leadZerosBin[1] ), 
         .Z(n330[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i8_3_lut.init = 16'hcaca;
    LUT4 i29386_4_lut (.A(n265), .B(n73795), .C(n70630), .D(\leadZerosBin[2] ), 
         .Z(n301[6])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i29386_4_lut.init = 16'h3022;
    LUT4 mux_26_i9_3_lut (.A(n301[8]), .B(n301[6]), .C(\leadZerosBin[1] ), 
         .Z(n330[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i9_3_lut.init = 16'hcaca;
    LUT4 mux_21_i10_3_lut (.A(n330[9]), .B(n330[8]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[9] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i10_3_lut.init = 16'hcaca;
    LUT4 mux_21_i9_3_lut (.A(n330[8]), .B(n330[7]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[8] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i9_3_lut.init = 16'hcaca;
    LUT4 i29575_4_lut (.A(\frac[7] ), .B(n70633), .C(n70707), .D(\leadZerosBin[2] ), 
         .Z(n301[7])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i29575_4_lut.init = 16'h3022;
    LUT4 mux_26_i10_3_lut (.A(n301[9]), .B(n301[7]), .C(\leadZerosBin[1] ), 
         .Z(n330[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i10_3_lut.init = 16'hcaca;
    LUT4 mux_26_i11_3_lut (.A(n301[10]), .B(n301[8]), .C(\leadZerosBin[1] ), 
         .Z(n330[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i11_3_lut.init = 16'hcaca;
    LUT4 mux_21_i12_3_lut (.A(n330[11]), .B(n330[10]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[11] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i12_3_lut.init = 16'hcaca;
    LUT4 mux_21_i11_3_lut (.A(n330[10]), .B(n330[9]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[10] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i11_3_lut.init = 16'hcaca;
    LUT4 mux_26_i12_3_lut (.A(n301[11]), .B(n301[9]), .C(\leadZerosBin[1] ), 
         .Z(n330[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i12_3_lut.init = 16'hcaca;
    LUT4 mux_26_i13_3_lut (.A(n301[12]), .B(n301[10]), .C(\leadZerosBin[1] ), 
         .Z(n330[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i13_3_lut.init = 16'hcaca;
    LUT4 mux_21_i14_3_lut (.A(n330[13]), .B(n330[12]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[13] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i14_3_lut.init = 16'hcaca;
    LUT4 mux_21_i13_3_lut (.A(n330[12]), .B(n330[11]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[12] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i13_3_lut.init = 16'hcaca;
    LUT4 mux_26_i14_4_lut (.A(n20408), .B(n301[11]), .C(\leadZerosBin[1] ), 
         .D(n70638), .Z(n330[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_26_i14_4_lut.init = 16'hcac0;
    LUT4 mux_30_i9_4_lut (.A(n263), .B(\addSubAB[0] ), .C(n73795), .D(n70637), 
         .Z(n272[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_30_i9_4_lut.init = 16'h0aca;
    LUT4 mux_28_i13_3_lut (.A(n272[12]), .B(n272[8]), .C(\leadZerosBin[2] ), 
         .Z(n301[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_28_i13_3_lut.init = 16'hcaca;
    LUT4 mux_26_i15_3_lut (.A(n301[14]), .B(n301[12]), .C(\leadZerosBin[1] ), 
         .Z(n330[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i15_3_lut.init = 16'hcaca;
    LUT4 mux_21_i16_3_lut (.A(n330[15]), .B(n330[14]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[15] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i16_3_lut.init = 16'hcaca;
    LUT4 mux_21_i15_3_lut (.A(n330[14]), .B(n330[13]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[14] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i15_3_lut.init = 16'hcaca;
    LUT4 i9067_3_lut (.A(n19134), .B(n19142), .C(\leadZerosBin[2] ), .Z(n20408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9067_3_lut.init = 16'hcaca;
    LUT4 i29635_4_lut (.A(n20404), .B(n70638), .C(n20408), .D(\leadZerosBin[1] ), 
         .Z(n330[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29635_4_lut.init = 16'hc088;
    LUT4 i29618_4_lut (.A(n19132), .B(n70638), .C(n19140), .D(\leadZerosBin[2] ), 
         .Z(n301[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29618_4_lut.init = 16'hc088;
    LUT4 mux_26_i17_3_lut (.A(n301[16]), .B(n301[14]), .C(\leadZerosBin[1] ), 
         .Z(n330[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i17_3_lut.init = 16'hcaca;
    LUT4 mux_21_i18_3_lut (.A(n330[17]), .B(n330[16]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i18_3_lut.init = 16'hcaca;
    LUT4 mux_21_i17_3_lut (.A(n330[16]), .B(n330[15]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i17_3_lut.init = 16'hcaca;
    LUT4 i9063_3_lut (.A(n19130), .B(n19138), .C(\leadZerosBin[2] ), .Z(n20404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9063_3_lut.init = 16'hcaca;
    LUT4 mux_26_i18_4_lut (.A(n301[17]), .B(n20404), .C(\leadZerosBin[1] ), 
         .D(n70638), .Z(n330[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_26_i18_4_lut.init = 16'hca0a;
    LUT4 i29391_4_lut (.A(\frac[12] ), .B(n70638), .C(n70706), .D(n73795), 
         .Z(n272[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29391_4_lut.init = 16'hc088;
    LUT4 mux_28_i17_3_lut (.A(n272[16]), .B(n272[12]), .C(\leadZerosBin[2] ), 
         .Z(n301[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_28_i17_3_lut.init = 16'hcaca;
    LUT4 mux_26_i19_3_lut (.A(n301[18]), .B(n301[16]), .C(\leadZerosBin[1] ), 
         .Z(n330[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i19_3_lut.init = 16'hcaca;
    LUT4 mux_21_i20_3_lut (.A(n330[19]), .B(n330[18]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[19] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i20_3_lut.init = 16'hcaca;
    LUT4 mux_21_i19_3_lut (.A(n330[18]), .B(n330[17]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[18] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i19_3_lut.init = 16'hcaca;
    LUT4 i7834_3_lut (.A(\frac[13] ), .B(n70703), .C(n73795), .Z(n19134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7834_3_lut.init = 16'hcaca;
    LUT4 mux_28_i18_4_lut (.A(n272[17]), .B(n19134), .C(\leadZerosBin[2] ), 
         .D(n70638), .Z(n301[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_28_i18_4_lut.init = 16'hca0a;
    LUT4 mux_26_i20_3_lut (.A(n301[19]), .B(n301[17]), .C(\leadZerosBin[1] ), 
         .Z(n330[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i20_3_lut.init = 16'hcaca;
    LUT4 i7832_3_lut (.A(\frac[14] ), .B(\frac[6] ), .C(n73795), .Z(n19132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7832_3_lut.init = 16'hcaca;
    LUT4 mux_28_i19_4_lut (.A(n272[18]), .B(n19132), .C(\leadZerosBin[2] ), 
         .D(n70638), .Z(n301[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_28_i19_4_lut.init = 16'hca0a;
    LUT4 mux_26_i21_3_lut (.A(n301[20]), .B(n301[18]), .C(\leadZerosBin[1] ), 
         .Z(n330[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i21_3_lut.init = 16'hcaca;
    LUT4 mux_21_i22_3_lut (.A(n330[21]), .B(n330[20]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i22_3_lut.init = 16'hcaca;
    LUT4 mux_21_i21_3_lut (.A(n330[20]), .B(n330[19]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[20] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i21_3_lut.init = 16'hcaca;
    LUT4 i7830_3_lut (.A(\frac[15] ), .B(\frac[7] ), .C(n73795), .Z(n19130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7830_3_lut.init = 16'hcaca;
    LUT4 mux_28_i20_4_lut (.A(n272[19]), .B(n19130), .C(\leadZerosBin[2] ), 
         .D(n70638), .Z(n301[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_28_i20_4_lut.init = 16'hca0a;
    LUT4 mux_26_i22_3_lut (.A(n301[21]), .B(n301[19]), .C(\leadZerosBin[1] ), 
         .Z(n330[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i22_3_lut.init = 16'hcaca;
    LUT4 mux_30_i17_3_lut (.A(n243[16]), .B(n263), .C(n73795), .Z(n272[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_30_i17_3_lut.init = 16'hcaca;
    LUT4 mux_28_i21_3_lut (.A(n272[20]), .B(n272[16]), .C(\leadZerosBin[2] ), 
         .Z(n301[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_28_i21_3_lut.init = 16'hcaca;
    LUT4 mux_26_i23_3_lut (.A(n301[22]), .B(n301[20]), .C(\leadZerosBin[1] ), 
         .Z(n330[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i23_3_lut.init = 16'hcaca;
    LUT4 mux_21_i24_3_lut (.A(n330[23]), .B(n330[22]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i24_3_lut.init = 16'hcaca;
    LUT4 mux_21_i23_3_lut (.A(n330[22]), .B(n330[21]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[22] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i23_3_lut.init = 16'hcaca;
    LUT4 mux_30_i18_4_lut (.A(n243[17]), .B(\frac[9] ), .C(n73795), .D(n70638), 
         .Z(n272[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam mux_30_i18_4_lut.init = 16'hca0a;
    LUT4 mux_28_i22_3_lut (.A(n272[21]), .B(n272[17]), .C(\leadZerosBin[2] ), 
         .Z(n301[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_28_i22_3_lut.init = 16'hcaca;
    LUT4 mux_26_i24_3_lut (.A(n301[23]), .B(n301[21]), .C(\leadZerosBin[1] ), 
         .Z(n330[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_26_i24_3_lut.init = 16'hcaca;
    LUT4 mux_21_i25_3_lut (.A(n330[24]), .B(n330[23]), .C(\leadZerosBin[0] ), 
         .Z(\frac_sub_Norm1[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_21_i25_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut_adj_758 (.A(n24_c), .B(n20), .C(n70674), .D(n18), 
         .Z(n62779)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_758.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_759 (.A(n66751), .B(n24_c), .C(n70685), .D(\frac[13] ), 
         .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_759.init = 16'hfffe;
    LUT4 i1_2_lut_rep_686_4_lut (.A(n66751), .B(n24_c), .C(n70685), .D(n23), 
         .Z(n70656)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_686_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_676_3_lut_4_lut (.A(n23), .B(n70662), .C(n70671), 
         .D(n27), .Z(n70646)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_676_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_28_i9_3_lut_4_lut (.A(n70706), .B(n70633), .C(\leadZerosBin[2] ), 
         .D(n272[8]), .Z(n301[8])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_28_i9_3_lut_4_lut.init = 16'h2f20;
    LUT4 i2_3_lut_4_lut_adj_760 (.A(n70650), .B(n70656), .C(n5), .D(n66650), 
         .Z(n66653)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_760.init = 16'h8000;
    LUT4 i30_3_lut_4_lut (.A(\leadZerosBin[1] ), .B(n70622), .C(\leadZerosBin[0] ), 
         .D(n19114), .Z(n17)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i30_3_lut_4_lut.init = 16'h4f40;
    LUT4 i1_3_lut_rep_673 (.A(n70703), .B(\frac[6] ), .C(n39), .Z(n70643)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_673.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_761 (.A(n70707), .B(n70706), .C(n70643), .D(n70714), 
         .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_761.init = 16'hfffe;
    LUT4 i1_3_lut_rep_671 (.A(n70707), .B(n70706), .C(n70643), .Z(n70641)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_671.init = 16'hfefe;
    LUT4 mux_53_i7_3_lut_else_3_lut (.A(\addSubAB[6] ), .B(\subBAExpEq[6] ), 
         .C(n70733), .Z(n70869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i7_3_lut_else_3_lut.init = 16'hcaca;
    LUT4 mux_53_i7_3_lut_then_3_lut (.A(\B_int[3] ), .B(\A_int[3] ), .C(n70737), 
         .Z(n70870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_53_i7_3_lut_then_3_lut.init = 16'hcaca;
    LUT4 i28179_2_lut_rep_693_4_lut (.A(\frac[20] ), .B(n66680), .C(\frac[21] ), 
         .D(n18), .Z(n70663)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i28179_2_lut_rep_693_4_lut.init = 16'heee0;
    LUT4 i1_2_lut_rep_698_3_lut (.A(\frac[19] ), .B(\frac[20] ), .C(n66680), 
         .Z(n70668)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_698_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\frac[19] ), .B(\frac[20] ), .C(n66680), 
         .D(n70672), .Z(n66650)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_704_4_lut (.A(\frac[25] ), .B(\frac[26] ), .C(\frac[23] ), 
         .D(\frac[24] ), .Z(n70674)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_704_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_715_4_lut (.A(\frac[18] ), .B(\frac[19] ), .C(\frac[16] ), 
         .D(\frac[17] ), .Z(n70685)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_715_4_lut.init = 16'hfffe;
    LUT4 mux_21_i3_3_lut_4_lut (.A(\leadZerosBin[2] ), .B(n70616), .C(\leadZerosBin[0] ), 
         .D(n356), .Z(\frac_sub_Norm1[2] )) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_21_i3_3_lut_4_lut.init = 16'h4f40;
    LUT4 i1_4_lut_4_lut_adj_762 (.A(\frac[25] ), .B(\frac[26] ), .C(\frac[23] ), 
         .D(\frac[24] ), .Z(n112)) /* synthesis lut_function=(!(A (B)+!A (B+((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_adj_762.init = 16'h2232;
    LUT4 n70128_bdd_2_lut_3_lut (.A(n70127), .B(\frac[8] ), .C(\frac[9] ), 
         .Z(n70129)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam n70128_bdd_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_3_lut (.A(\frac[9] ), .B(\frac[10] ), .C(n31), .Z(n35)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_763 (.A(\frac[7] ), .B(\frac[8] ), .C(\frac[9] ), 
         .D(n22464), .Z(n39)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_763.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module \right_shifter(27,8,4)_U27 
//

module \right_shifter(27,8,4)_U27  (diffExpAB, diffExpBA, \diffExp[4] , 
            n70777, n70835, \B_int[19] , \A_int[19] , n70834, \B_int[15] , 
            \A_int[15] , n70833, n70832, \B_int[1] , \A_int[1] , \diffExp[2] , 
            \efectFracB[21] , \efectFracB[20] , n70743, \efectFracB[19] , 
            \efectFracB[15] , \efectFracB[16] , n19214, n15, n28, 
            n66904, n70771, n9, \efectFracB[14] , \efectFracB[7] , 
            \efectFracB[5] , \efectFracB[12] , n70820, \efectFracB[13] , 
            n27, \fracAlign_int[0] , n70740, n7, \efectFracB_align[2] , 
            \efectFracB_align[1] , \B_int[0] , \A_int[0] , \fracAlign_int[4] , 
            \fracAlign_int[3] , n55, \fracAlign_int[6] , \fracAlign_int[5] , 
            \B_int[5] , \A_int[5] , \fracAlign_int[8] , \fracAlign_int[7] , 
            \B_int[6] , \A_int[6] , \fracAlign_int[10] , \fracAlign_int[9] , 
            \B_int[8] , \A_int[8] , \fracAlign_int[12] , n41778, \fracAlign_int[14] , 
            \fracAlign_int[13] , \fracAlign_int[16] , \fracAlign_int[15] , 
            \fracAlign_int[18] , \fracAlign_int[17] , \fracAlign_int[20] , 
            n41588, \fracAlign_int[22] , \fracAlign_int[21] , n66914, 
            n66178, \B_int[22] , \A_int[22] , \B_int[14] , \A_int[14] , 
            \B_int[21] , \A_int[21] , \B_int[20] , \A_int[20] );
    input [8:0]diffExpAB;
    input [8:0]diffExpBA;
    output \diffExp[4] ;
    output n70777;
    output n70835;
    input \B_int[19] ;
    input \A_int[19] ;
    output n70834;
    input \B_int[15] ;
    input \A_int[15] ;
    output n70833;
    output n70832;
    input \B_int[1] ;
    input \A_int[1] ;
    output \diffExp[2] ;
    input \efectFracB[21] ;
    input \efectFracB[20] ;
    output n70743;
    input \efectFracB[19] ;
    input \efectFracB[15] ;
    input \efectFracB[16] ;
    input n19214;
    output n15;
    input n28;
    output n66904;
    input n70771;
    input n9;
    input \efectFracB[14] ;
    input \efectFracB[7] ;
    input \efectFracB[5] ;
    input \efectFracB[12] ;
    input n70820;
    input \efectFracB[13] ;
    input n27;
    output \fracAlign_int[0] ;
    input n70740;
    output n7;
    output \efectFracB_align[2] ;
    output \efectFracB_align[1] ;
    input \B_int[0] ;
    input \A_int[0] ;
    output \fracAlign_int[4] ;
    output \fracAlign_int[3] ;
    input n55;
    output \fracAlign_int[6] ;
    output \fracAlign_int[5] ;
    input \B_int[5] ;
    input \A_int[5] ;
    output \fracAlign_int[8] ;
    output \fracAlign_int[7] ;
    input \B_int[6] ;
    input \A_int[6] ;
    output \fracAlign_int[10] ;
    output \fracAlign_int[9] ;
    input \B_int[8] ;
    input \A_int[8] ;
    output \fracAlign_int[12] ;
    output n41778;
    output \fracAlign_int[14] ;
    output \fracAlign_int[13] ;
    output \fracAlign_int[16] ;
    output \fracAlign_int[15] ;
    output \fracAlign_int[18] ;
    output \fracAlign_int[17] ;
    output \fracAlign_int[20] ;
    output n41588;
    output \fracAlign_int[22] ;
    output \fracAlign_int[21] ;
    output n66914;
    output n66178;
    input \B_int[22] ;
    input \A_int[22] ;
    input \B_int[14] ;
    input \A_int[14] ;
    input \B_int[21] ;
    input \A_int[21] ;
    input \B_int[20] ;
    input \A_int[20] ;
    
    wire [27:0]efectFracB;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(67[23:33])
    wire [8:0]diffExp;   // c:/users/yisong/documents/new/mlp/fp_add.vhd(68[33:40])
    
    wire n70770, n70772, n14, n70819;
    wire [27:0]n69;
    wire [27:0]n37;
    
    wire n66626, n70776, n70775, n70774, n41656, n70773, n20420, 
        n41436;
    wire [27:0]n5;
    
    wire n11, n6;
    wire [27:0]n101;
    
    wire n9_c, n19865, n66931, n66933, n22, n21, n23, n63170, 
        n66999, n34, n19218, n19220, n19216, n20428, n20426, n20606, 
        n20424, n41736, n20422, n20604, n23579, n70923, n70924;
    
    LUT4 i28411_2_lut_rep_807_4_lut (.A(diffExpAB[3]), .B(diffExpBA[3]), 
         .C(diffExpAB[8]), .D(\diffExp[4] ), .Z(n70777)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i28411_2_lut_rep_807_4_lut.init = 16'hffca;
    LUT4 mux_2997_i4_3_lut_rep_865 (.A(diffExpAB[3]), .B(diffExpBA[3]), 
         .C(diffExpAB[8]), .Z(n70835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2997_i4_3_lut_rep_865.init = 16'hcaca;
    LUT4 mux_3876_i20_3_lut_rep_864 (.A(\B_int[19] ), .B(\A_int[19] ), .C(diffExpAB[8]), 
         .Z(n70834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i20_3_lut_rep_864.init = 16'hcaca;
    LUT4 i28281_2_lut_rep_800_4_lut (.A(\B_int[15] ), .B(\A_int[15] ), .C(diffExpAB[8]), 
         .D(\diffExp[4] ), .Z(n70770)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i28281_2_lut_rep_800_4_lut.init = 16'hca00;
    LUT4 mux_3876_i16_3_lut_rep_863 (.A(\B_int[15] ), .B(\A_int[15] ), .C(diffExpAB[8]), 
         .Z(n70833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i16_3_lut_rep_863.init = 16'hcaca;
    LUT4 i1_2_lut_rep_802_4_lut (.A(diffExpAB[1]), .B(diffExpBA[1]), .C(diffExpAB[8]), 
         .D(efectFracB[24]), .Z(n70772)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_802_4_lut.init = 16'hffca;
    LUT4 mux_2997_i2_3_lut_rep_862 (.A(diffExpAB[1]), .B(diffExpBA[1]), 
         .C(diffExpAB[8]), .Z(n70832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2997_i2_3_lut_rep_862.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(\B_int[1] ), .B(\A_int[1] ), .C(diffExpAB[8]), 
         .D(efectFracB[11]), .Z(n14)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_3876_i2_3_lut_rep_849 (.A(\B_int[1] ), .B(\A_int[1] ), .C(diffExpAB[8]), 
         .Z(n70819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i2_3_lut_rep_849.init = 16'hcaca;
    LUT4 i29585_2_lut_3_lut_4_lut (.A(\diffExp[4] ), .B(n70835), .C(efectFracB[24]), 
         .D(\diffExp[2] ), .Z(n69[24])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i29585_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i29586_2_lut_3_lut_4_lut (.A(\diffExp[4] ), .B(n70835), .C(efectFracB[23]), 
         .D(\diffExp[2] ), .Z(n69[23])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i29586_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut (.A(\diffExp[4] ), .B(n70835), .C(\efectFracB[21] ), 
         .Z(n37[21])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_736 (.A(\diffExp[4] ), .B(n70835), .C(\efectFracB[20] ), 
         .Z(n37[20])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_736.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\diffExp[4] ), .B(n70835), .C(n70834), 
         .D(\diffExp[2] ), .Z(n66626)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i53877_2_lut_rep_773_3_lut (.A(\diffExp[4] ), .B(n70835), .C(\diffExp[2] ), 
         .Z(n70743)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i53877_2_lut_rep_773_3_lut.init = 16'hfefe;
    LUT4 i29410_2_lut_3_lut (.A(\diffExp[4] ), .B(n70835), .C(\efectFracB[19] ), 
         .Z(n37[19])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29410_2_lut_3_lut.init = 16'h1010;
    LUT4 i29409_2_lut_3_lut (.A(\diffExp[4] ), .B(n70835), .C(n70834), 
         .Z(n37[22])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29409_2_lut_3_lut.init = 16'h1010;
    LUT4 i29413_2_lut_4_lut (.A(\efectFracB[15] ), .B(efectFracB[23]), .C(n70835), 
         .D(\diffExp[4] ), .Z(n37[15])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29413_2_lut_4_lut.init = 16'h00ca;
    LUT4 i7912_3_lut_rep_806 (.A(\efectFracB[15] ), .B(efectFracB[23]), 
         .C(n70835), .Z(n70776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7912_3_lut_rep_806.init = 16'hcaca;
    LUT4 i29412_2_lut_4_lut (.A(\efectFracB[16] ), .B(efectFracB[24]), .C(n70835), 
         .D(\diffExp[4] ), .Z(n37[16])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29412_2_lut_4_lut.init = 16'h00ca;
    LUT4 i7910_3_lut_rep_805 (.A(\efectFracB[16] ), .B(efectFracB[24]), 
         .C(n70835), .Z(n70775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7910_3_lut_rep_805.init = 16'hcaca;
    LUT4 i29411_2_lut_4_lut (.A(efectFracB[17]), .B(efectFracB[25]), .C(n70835), 
         .D(\diffExp[4] ), .Z(n37[17])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29411_2_lut_4_lut.init = 16'h00ca;
    LUT4 i7908_3_lut_rep_804 (.A(efectFracB[17]), .B(efectFracB[25]), .C(n70835), 
         .Z(n70774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7908_3_lut_rep_804.init = 16'hcaca;
    LUT4 mux_3900_i15_3_lut_4_lut (.A(n70835), .B(n70833), .C(\diffExp[2] ), 
         .D(n19214), .Z(n41656)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3900_i15_3_lut_4_lut.init = 16'hefe0;
    LUT4 i29844_2_lut_3_lut (.A(n70835), .B(n70833), .C(\diffExp[4] ), 
         .Z(n37[18])) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i29844_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i29630_2_lut_4_lut (.A(\efectFracB[21] ), .B(efectFracB[25]), .C(\diffExp[2] ), 
         .D(n70777), .Z(n69[21])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i29630_2_lut_4_lut.init = 16'h00ca;
    LUT4 i9077_3_lut_rep_803 (.A(\efectFracB[21] ), .B(efectFracB[25]), 
         .C(\diffExp[2] ), .Z(n70773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9077_3_lut_rep_803.init = 16'hcaca;
    LUT4 i9073_3_lut_4_lut (.A(\diffExp[2] ), .B(n70834), .C(n70832), 
         .D(n20420), .Z(n41436)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i9073_3_lut_4_lut.init = 16'hefe0;
    LUT4 i24_4_lut_4_lut (.A(efectFracB[24]), .B(n70832), .C(diffExp[0]), 
         .D(efectFracB[25]), .Z(n15)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam i24_4_lut_4_lut.init = 16'h3e0e;
    LUT4 i4_3_lut_4_lut (.A(n70833), .B(\diffExp[4] ), .C(n5[7]), .D(n28), 
         .Z(n11)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i4_3_lut_4_lut.init = 16'hfff8;
    LUT4 i53998_3_lut_4_lut (.A(\diffExp[2] ), .B(n70777), .C(efectFracB[25]), 
         .D(diffExp[0]), .Z(n66904)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i53998_3_lut_4_lut.init = 16'h1110;
    LUT4 i2_2_lut_4_lut (.A(n70770), .B(n70771), .C(n70835), .D(n37[3]), 
         .Z(n6)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i2_2_lut_4_lut.init = 16'hffca;
    PFUMX mux_3900_i16 (.BLUT(n37[15]), .ALUT(n37[19]), .C0(\diffExp[2] ), 
          .Z(n69[15]));
    PFUMX mux_3900_i17 (.BLUT(n37[16]), .ALUT(n37[20]), .C0(\diffExp[2] ), 
          .Z(n69[16]));
    PFUMX mux_3900_i18 (.BLUT(n37[17]), .ALUT(n37[21]), .C0(\diffExp[2] ), 
          .Z(n69[17]));
    PFUMX mux_3900_i19 (.BLUT(n37[18]), .ALUT(n37[22]), .C0(\diffExp[2] ), 
          .Z(n69[18]));
    PFUMX mux_3905_i22 (.BLUT(n69[21]), .ALUT(n69[23]), .C0(n70832), .Z(n101[21]));
    PFUMX mux_3905_i23 (.BLUT(n66626), .ALUT(n69[24]), .C0(n70832), .Z(n101[22]));
    LUT4 mux_3900_i1_3_lut (.A(n37[0]), .B(n37[4]), .C(\diffExp[2] ), 
         .Z(n69[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i1_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i1_4_lut (.A(\diffExp[4] ), .B(n5[8]), .C(n70835), .D(\efectFracB[16] ), 
         .Z(n37[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3895_i1_4_lut.init = 16'hcac0;
    LUT4 i2_4_lut (.A(\diffExp[4] ), .B(n5[3]), .C(efectFracB[17]), .D(\efectFracB[16] ), 
         .Z(n9_c)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i2_4_lut.init = 16'heeec;
    LUT4 i8563_4_lut (.A(\diffExp[2] ), .B(n37[0]), .C(n6), .D(n37[1]), 
         .Z(n19865)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i8563_4_lut.init = 16'haaa8;
    LUT4 i54023_3_lut (.A(n70832), .B(n69[0]), .C(n69[1]), .Z(n66931)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i54023_3_lut.init = 16'ha8a8;
    LUT4 i54025_4_lut (.A(n69[0]), .B(n19865), .C(n69[2]), .D(n70832), 
         .Z(n66933)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i54025_4_lut.init = 16'hfcee;
    LUT4 i9_4_lut (.A(n9), .B(\efectFracB[14] ), .C(efectFracB[3]), .D(\efectFracB[7] ), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(\efectFracB[15] ), .B(\efectFracB[5] ), .C(efectFracB[8]), 
         .D(\efectFracB[12] ), .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(n70820), .B(\efectFracB[13] ), .C(efectFracB[9]), 
         .D(n14), .Z(n23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(n11), .B(n9_c), .C(n27), .D(n5[4]), .Z(n63170)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i54090_4_lut (.A(n101[1]), .B(n66933), .C(n66931), .D(diffExp[0]), 
         .Z(n66999)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i54090_4_lut.init = 16'hfefc;
    LUT4 i27809_4_lut (.A(n23), .B(\diffExp[4] ), .C(n21), .D(n22), 
         .Z(n34)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i27809_4_lut.init = 16'hccc8;
    LUT4 i54112_4_lut (.A(n34), .B(n66999), .C(n63170), .D(n70835), 
         .Z(\fracAlign_int[0] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i54112_4_lut.init = 16'hfeee;
    LUT4 mux_3900_i3_3_lut (.A(n70740), .B(n37[6]), .C(\diffExp[2] ), 
         .Z(n69[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i3_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i2_4_lut (.A(\diffExp[4] ), .B(n5[9]), .C(n70835), .D(efectFracB[17]), 
         .Z(n37[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_3895_i2_4_lut.init = 16'hcac0;
    LUT4 mux_3900_i2_3_lut (.A(n37[1]), .B(n37[5]), .C(\diffExp[2] ), 
         .Z(n69[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i2_3_lut (.A(n69[1]), .B(n69[3]), .C(n70832), .Z(n101[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i3_3_lut (.A(n69[2]), .B(n69[4]), .C(n70832), .Z(n101[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i3_3_lut.init = 16'hcaca;
    LUT4 i28274_4_lut (.A(n101[2]), .B(n7), .C(n101[3]), .D(diffExp[0]), 
         .Z(\efectFracB_align[2] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i28274_4_lut.init = 16'h3022;
    LUT4 i28275_4_lut (.A(n101[1]), .B(n7), .C(n101[2]), .D(diffExp[0]), 
         .Z(\efectFracB_align[1] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i28275_4_lut.init = 16'h3022;
    LUT4 mux_3876_i1_3_lut (.A(\B_int[0] ), .B(\A_int[0] ), .C(diffExpAB[8]), 
         .Z(efectFracB[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i1_3_lut.init = 16'hcaca;
    LUT4 mux_3890_i4_3_lut (.A(efectFracB[3]), .B(\efectFracB[19] ), .C(\diffExp[4] ), 
         .Z(n5[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3890_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i4_4_lut (.A(n5[3]), .B(efectFracB[11]), .C(n70835), 
         .D(\diffExp[4] ), .Z(n37[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3895_i4_4_lut.init = 16'h0aca;
    LUT4 mux_3900_i4_3_lut (.A(n37[3]), .B(n37[7]), .C(\diffExp[2] ), 
         .Z(n69[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i4_3_lut (.A(n69[3]), .B(n69[5]), .C(n70832), .Z(n101[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3890_i5_3_lut (.A(n70819), .B(\efectFracB[20] ), .C(\diffExp[4] ), 
         .Z(n5[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3890_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i5_4_lut (.A(n5[4]), .B(\diffExp[4] ), .C(n70835), .D(\efectFracB[12] ), 
         .Z(n37[4])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3895_i5_4_lut.init = 16'h3a0a;
    LUT4 mux_3900_i5_3_lut (.A(n37[4]), .B(n37[8]), .C(\diffExp[2] ), 
         .Z(n69[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i5_3_lut (.A(n69[4]), .B(n69[6]), .C(n70832), .Z(n101[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i5_3_lut (.A(n101[4]), .B(n101[5]), .C(diffExp[0]), 
         .Z(\fracAlign_int[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i4_3_lut (.A(n101[3]), .B(n101[4]), .C(diffExp[0]), 
         .Z(\fracAlign_int[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i7_4_lut (.A(n27), .B(\diffExp[4] ), .C(n70835), .D(\efectFracB[14] ), 
         .Z(n37[6])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3895_i7_4_lut.init = 16'h3a0a;
    LUT4 mux_3900_i7_3_lut (.A(n37[6]), .B(n55), .C(\diffExp[2] ), .Z(n69[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i6_4_lut (.A(n28), .B(\diffExp[4] ), .C(n70835), .D(\efectFracB[13] ), 
         .Z(n37[5])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3895_i6_4_lut.init = 16'h3a0a;
    LUT4 mux_3900_i6_3_lut (.A(n37[5]), .B(n37[9]), .C(\diffExp[2] ), 
         .Z(n69[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3900_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i6_3_lut (.A(n69[5]), .B(n69[7]), .C(n70832), .Z(n101[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i7_3_lut (.A(n69[6]), .B(n69[8]), .C(n70832), .Z(n101[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i7_3_lut (.A(n101[6]), .B(n101[7]), .C(diffExp[0]), 
         .Z(\fracAlign_int[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i6_3_lut (.A(n101[5]), .B(n101[6]), .C(diffExp[0]), 
         .Z(\fracAlign_int[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3876_i6_3_lut (.A(\B_int[5] ), .B(\A_int[5] ), .C(diffExpAB[8]), 
         .Z(efectFracB[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3890_i9_3_lut (.A(efectFracB[8]), .B(efectFracB[24]), .C(\diffExp[4] ), 
         .Z(n5[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3890_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i9_4_lut (.A(n5[8]), .B(\diffExp[4] ), .C(n70835), .D(\efectFracB[16] ), 
         .Z(n37[8])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3895_i9_4_lut.init = 16'h3a0a;
    LUT4 mux_3900_i9_4_lut (.A(n37[8]), .B(n19218), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3900_i9_4_lut.init = 16'h0aca;
    LUT4 mux_3890_i8_3_lut (.A(\efectFracB[7] ), .B(efectFracB[23]), .C(\diffExp[4] ), 
         .Z(n5[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3890_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i8_4_lut (.A(n5[7]), .B(\diffExp[4] ), .C(n70835), .D(\efectFracB[15] ), 
         .Z(n37[7])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3895_i8_4_lut.init = 16'h3a0a;
    LUT4 mux_3900_i8_4_lut (.A(n37[7]), .B(n19220), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3900_i8_4_lut.init = 16'h0aca;
    LUT4 mux_3905_i8_3_lut (.A(n69[7]), .B(n69[9]), .C(n70832), .Z(n101[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i9_3_lut (.A(n69[8]), .B(n69[10]), .C(n70832), .Z(n101[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i9_3_lut (.A(n101[8]), .B(n101[9]), .C(diffExp[0]), 
         .Z(\fracAlign_int[8] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i9_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i8_3_lut (.A(n101[7]), .B(n101[8]), .C(diffExp[0]), 
         .Z(\fracAlign_int[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3900_i11_4_lut (.A(n55), .B(n19214), .C(\diffExp[2] ), .D(\diffExp[4] ), 
         .Z(n69[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3900_i11_4_lut.init = 16'h0aca;
    LUT4 mux_3876_i7_3_lut (.A(\B_int[6] ), .B(\A_int[6] ), .C(diffExpAB[8]), 
         .Z(efectFracB[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3890_i10_3_lut (.A(efectFracB[9]), .B(efectFracB[25]), .C(\diffExp[4] ), 
         .Z(n5[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3890_i10_3_lut.init = 16'hcaca;
    LUT4 mux_3895_i10_4_lut (.A(n5[9]), .B(\diffExp[4] ), .C(n70835), 
         .D(efectFracB[17]), .Z(n37[9])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam mux_3895_i10_4_lut.init = 16'h3a0a;
    LUT4 mux_3900_i10_4_lut (.A(n37[9]), .B(n19216), .C(\diffExp[2] ), 
         .D(\diffExp[4] ), .Z(n69[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3900_i10_4_lut.init = 16'h0aca;
    LUT4 mux_3905_i10_4_lut (.A(n69[9]), .B(n20428), .C(n70832), .D(\diffExp[4] ), 
         .Z(n101[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3905_i10_4_lut.init = 16'h0aca;
    LUT4 mux_3905_i11_4_lut (.A(n69[10]), .B(n20426), .C(n70832), .D(\diffExp[4] ), 
         .Z(n101[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3905_i11_4_lut.init = 16'h0aca;
    LUT4 mux_3910_i11_4_lut (.A(n101[10]), .B(n20606), .C(diffExp[0]), 
         .D(\diffExp[4] ), .Z(\fracAlign_int[10] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3910_i11_4_lut.init = 16'h0aca;
    LUT4 mux_3910_i10_3_lut (.A(n101[9]), .B(n101[10]), .C(diffExp[0]), 
         .Z(\fracAlign_int[9] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i10_3_lut.init = 16'hcaca;
    LUT4 i7918_3_lut (.A(\efectFracB[12] ), .B(\efectFracB[20] ), .C(n70835), 
         .Z(n19218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7918_3_lut.init = 16'hcaca;
    LUT4 i9085_3_lut (.A(n19218), .B(n70775), .C(\diffExp[2] ), .Z(n20426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9085_3_lut.init = 16'hcaca;
    LUT4 mux_3876_i9_3_lut (.A(\B_int[8] ), .B(\A_int[8] ), .C(diffExpAB[8]), 
         .Z(efectFracB[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i9_3_lut.init = 16'hcaca;
    LUT4 i7920_3_lut (.A(efectFracB[11]), .B(\efectFracB[19] ), .C(n70835), 
         .Z(n19220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7920_3_lut.init = 16'hcaca;
    LUT4 i9087_3_lut (.A(n19220), .B(n70776), .C(\diffExp[2] ), .Z(n20428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9087_3_lut.init = 16'hcaca;
    LUT4 i9261_3_lut (.A(n20428), .B(n20424), .C(n70832), .Z(n20606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9261_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i13_3_lut (.A(n20426), .B(n41656), .C(n70832), .Z(n41736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i13_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i13_4_lut (.A(\diffExp[4] ), .B(n101[13]), .C(diffExp[0]), 
         .D(n41736), .Z(\fracAlign_int[12] )) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3910_i13_4_lut.init = 16'hc5c0;
    LUT4 mux_3910_i12_3_lut (.A(n20606), .B(n41736), .C(diffExp[0]), .Z(n41778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i12_3_lut.init = 16'hcaca;
    LUT4 i7916_3_lut (.A(\efectFracB[13] ), .B(\efectFracB[21] ), .C(n70835), 
         .Z(n19216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7916_3_lut.init = 16'hcaca;
    LUT4 i9083_3_lut (.A(n19216), .B(n70774), .C(\diffExp[2] ), .Z(n20424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9083_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i14_4_lut (.A(n20424), .B(n69[15]), .C(n70832), .D(\diffExp[4] ), 
         .Z(n101[13])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam mux_3905_i14_4_lut.init = 16'hc0ca;
    LUT4 mux_3905_i15_4_lut (.A(\diffExp[4] ), .B(n69[16]), .C(n70832), 
         .D(n41656), .Z(n101[14])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3905_i15_4_lut.init = 16'hc5c0;
    LUT4 mux_3910_i15_3_lut (.A(n101[14]), .B(n101[15]), .C(diffExp[0]), 
         .Z(\fracAlign_int[14] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i15_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i14_3_lut (.A(n101[13]), .B(n101[14]), .C(diffExp[0]), 
         .Z(\fracAlign_int[13] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i14_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i16_3_lut (.A(n69[15]), .B(n69[17]), .C(n70832), .Z(n101[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i16_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i17_3_lut (.A(n69[16]), .B(n69[18]), .C(n70832), .Z(n101[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3905_i17_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i17_3_lut (.A(n101[16]), .B(n101[17]), .C(diffExp[0]), 
         .Z(\fracAlign_int[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i17_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i16_3_lut (.A(n101[15]), .B(n101[16]), .C(diffExp[0]), 
         .Z(\fracAlign_int[15] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i16_3_lut.init = 16'hcaca;
    LUT4 mux_3905_i18_4_lut (.A(n69[17]), .B(n20422), .C(n70832), .D(n70777), 
         .Z(n101[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3905_i18_4_lut.init = 16'h0aca;
    LUT4 mux_3905_i19_4_lut (.A(n69[18]), .B(n20420), .C(n70832), .D(n70777), 
         .Z(n101[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3905_i19_4_lut.init = 16'h0aca;
    LUT4 mux_3910_i19_4_lut (.A(n101[18]), .B(n20604), .C(diffExp[0]), 
         .D(n70777), .Z(\fracAlign_int[18] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3910_i19_4_lut.init = 16'h0aca;
    LUT4 mux_3910_i18_3_lut (.A(n101[17]), .B(n101[18]), .C(diffExp[0]), 
         .Z(\fracAlign_int[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i18_3_lut.init = 16'hcaca;
    LUT4 i9079_3_lut (.A(\efectFracB[20] ), .B(efectFracB[24]), .C(\diffExp[2] ), 
         .Z(n20420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9079_3_lut.init = 16'hcaca;
    LUT4 i9081_3_lut (.A(\efectFracB[19] ), .B(efectFracB[23]), .C(\diffExp[2] ), 
         .Z(n20422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9081_3_lut.init = 16'hcaca;
    LUT4 i9259_3_lut (.A(n20422), .B(n70773), .C(n70832), .Z(n20604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9259_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i21_4_lut (.A(n41436), .B(n101[21]), .C(diffExp[0]), 
         .D(n70777), .Z(\fracAlign_int[20] )) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam mux_3910_i21_4_lut.init = 16'hc0ca;
    LUT4 i9257_3_lut (.A(n20604), .B(n41436), .C(diffExp[0]), .Z(n41588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i9257_3_lut.init = 16'hcaca;
    LUT4 mux_3910_i23_4_lut (.A(n101[22]), .B(n23579), .C(diffExp[0]), 
         .D(n70743), .Z(\fracAlign_int[22] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_3910_i23_4_lut.init = 16'h0aca;
    LUT4 mux_3910_i22_3_lut (.A(n101[21]), .B(n101[22]), .C(diffExp[0]), 
         .Z(\fracAlign_int[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3910_i22_3_lut.init = 16'hcaca;
    LUT4 i11896_3_lut (.A(efectFracB[23]), .B(efectFracB[25]), .C(n70832), 
         .Z(n23579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11896_3_lut.init = 16'hcaca;
    LUT4 i54006_4_lut (.A(n70777), .B(n23579), .C(n70772), .D(diffExp[0]), 
         .Z(n66914)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i54006_4_lut.init = 16'h5044;
    LUT4 mux_2997_i1_3_lut (.A(diffExpAB[0]), .B(diffExpBA[0]), .C(diffExpAB[8]), 
         .Z(diffExp[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2997_i1_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(n7), .B(n70743), .C(diffExp[0]), .D(n70832), .Z(n66178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    PFUMX i56112 (.BLUT(n70923), .ALUT(n70924), .C0(diffExpAB[8]), .Z(n7));
    LUT4 i3_4_lut_else_4_lut (.A(diffExpAB[5]), .B(diffExpAB[7]), .C(diffExpAB[6]), 
         .Z(n70923)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_4_lut_else_4_lut.init = 16'hfefe;
    LUT4 i3_4_lut_then_4_lut (.A(diffExpBA[7]), .B(diffExpBA[8]), .C(diffExpBA[6]), 
         .D(diffExpBA[5]), .Z(n70924)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_then_4_lut.init = 16'hfffe;
    LUT4 mux_3876_i23_3_lut (.A(\B_int[22] ), .B(\A_int[22] ), .C(diffExpAB[8]), 
         .Z(efectFracB[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i23_3_lut.init = 16'hcaca;
    LUT4 mux_3876_i15_3_lut (.A(\B_int[14] ), .B(\A_int[14] ), .C(diffExpAB[8]), 
         .Z(efectFracB[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i15_3_lut.init = 16'hcaca;
    LUT4 mux_3876_i22_3_lut (.A(\B_int[21] ), .B(\A_int[21] ), .C(diffExpAB[8]), 
         .Z(efectFracB[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i22_3_lut.init = 16'hcaca;
    LUT4 mux_3876_i21_3_lut (.A(\B_int[20] ), .B(\A_int[20] ), .C(diffExpAB[8]), 
         .Z(efectFracB[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_3876_i21_3_lut.init = 16'hcaca;
    LUT4 mux_2997_i5_3_lut (.A(diffExpAB[4]), .B(diffExpBA[4]), .C(diffExpAB[8]), 
         .Z(\diffExp[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2997_i5_3_lut.init = 16'hcaca;
    LUT4 mux_2997_i3_3_lut (.A(diffExpAB[2]), .B(diffExpBA[2]), .C(diffExpAB[8]), 
         .Z(\diffExp[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2997_i3_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module test
//

module test (sram_address_B, clock, GND_net, sram_output_B, n4599, 
            float_alu_c, i, n15113, n4617, n14054, n70822, \mlp_outputs[0] , 
            \mlp_outputs[1] , n23653, SDA_c, sram_ready_B, n23655, 
            weight_done, n2086, n70866, float_alu_ready, float_alu_b, 
            n927, n926, n70778, n70788, n14050, n2889, n3044, 
            n236, n61382, n63111, n23661, \float_alu_mode[1] , n27939, 
            n63112, \i[8] , \i[9] , n929, n928, \buf_r[83] , \buf_x[83] , 
            n2082, n73818, n923, n922, \state[0] , \float_alu_mode[2] , 
            n1155, n124, n2036, n70816, n2050, n2072, n2084, \i[12] , 
            \i[11] , \i[7] , \i[6] , \i[5] , \i[4] , \i[3] , n70716, 
            n24013, n62900, n932, n930, n63130, \buf_r[84] , \buf_x[84] , 
            \buf_r[85] , \buf_x[85] , \buf_r[86] , \buf_x[86] , \buf_r[87] , 
            \buf_x[87] , \buf_r[88] , \buf_x[88] , \buf_r[89] , \buf_x[89] , 
            n63113, mlp_done, n73801, n3946, n3944, n22106, n3961, 
            n62966, n62964, n63150, n63147, n63139, n63131, n63128, 
            n63122, n63120, n63116, n63115, n63109, n63114, n63107, 
            n63105, n63106, n63104, n63103, n63102, n62961, n63070, 
            n63069, n63156, n66524, n66522, n62958, n63068, n70867, 
            n921, n23942, n3988, n28181, n66628, n23639, n1156, 
            n73809, n45598, n931, n925, n924);
    output [11:0]sram_address_B;
    input clock;
    input GND_net;
    input [31:0]sram_output_B;
    input n4599;
    input [31:0]float_alu_c;
    output [31:0]i;
    input n15113;
    input n4617;
    output n14054;
    input n70822;
    output [31:0]\mlp_outputs[0] ;
    output [31:0]\mlp_outputs[1] ;
    input n23653;
    input SDA_c;
    output sram_ready_B;
    input n23655;
    input weight_done;
    output n2086;
    input n70866;
    output float_alu_ready;
    output [31:0]float_alu_b;
    input n927;
    input n926;
    input n70778;
    input n70788;
    output n14050;
    input [4:0]n2889;
    input [4:0]n3044;
    input [3:0]n236;
    input n61382;
    output n63111;
    output n23661;
    output \float_alu_mode[1] ;
    output n27939;
    output n63112;
    output \i[8] ;
    output \i[9] ;
    input n929;
    input n928;
    output \buf_r[83] ;
    input \buf_x[83] ;
    output n2082;
    input n73818;
    input n923;
    input n922;
    input \state[0] ;
    output \float_alu_mode[2] ;
    input n1155;
    output n124;
    output n2036;
    input n70816;
    output n2050;
    output n2072;
    output n2084;
    output \i[12] ;
    output \i[11] ;
    output \i[7] ;
    output \i[6] ;
    output \i[5] ;
    output \i[4] ;
    output \i[3] ;
    output n70716;
    output n24013;
    output n62900;
    input n932;
    input n930;
    output n63130;
    output \buf_r[84] ;
    input \buf_x[84] ;
    output \buf_r[85] ;
    input \buf_x[85] ;
    output \buf_r[86] ;
    input \buf_x[86] ;
    output \buf_r[87] ;
    input \buf_x[87] ;
    output \buf_r[88] ;
    input \buf_x[88] ;
    output \buf_r[89] ;
    input \buf_x[89] ;
    output n63113;
    output mlp_done;
    input n73801;
    input n3946;
    input n3944;
    output n22106;
    output n3961;
    output n62966;
    output n62964;
    output n63150;
    output n63147;
    output n63139;
    output n63131;
    output n63128;
    output n63122;
    output n63120;
    output n63116;
    output n63115;
    output n63109;
    output n63114;
    output n63107;
    output n63105;
    output n63106;
    output n63104;
    output n63103;
    output n63102;
    output n62961;
    output n63070;
    output n63069;
    output n63156;
    output n66524;
    output n66522;
    output n62958;
    output n63068;
    output n70867;
    input n921;
    output n23942;
    input n3988;
    input n28181;
    output n66628;
    output n23639;
    input n1156;
    input n73809;
    output n45598;
    input n931;
    input n925;
    input n924;
    
    wire [31:0]\temp_outputs[1] ;   // c:/users/yisong/documents/new/mlp/test.vhd(92[8:20])
    wire [31:0]\hidden_outputs[1] ;   // c:/users/yisong/documents/new/mlp/test.vhd(91[8:22])
    wire [31:0]h;   // c:/users/yisong/documents/new/mlp/test.vhd(166[11:12])
    wire [31:0]n;   // c:/users/yisong/documents/new/mlp/test.vhd(166[17:18])
    wire [31:0]\temp_outputs[0] ;   // c:/users/yisong/documents/new/mlp/test.vhd(92[8:20])
    wire [31:0]\hidden_outputs[0] ;   // c:/users/yisong/documents/new/mlp/test.vhd(91[8:22])
    wire [31:0]weight;   // c:/users/yisong/documents/new/mlp/test.vhd(172[8:14])
    wire [31:0]e;   // c:/users/yisong/documents/new/mlp/test.vhd(171[11:12])
    wire [31:0]addr;   // c:/users/yisong/documents/new/mlp/test.vhd(173[8:12])
    wire [31:0]\temp_outputs[4] ;   // c:/users/yisong/documents/new/mlp/test.vhd(92[8:20])
    wire [31:0]\hidden_outputs[4] ;   // c:/users/yisong/documents/new/mlp/test.vhd(91[8:22])
    wire [31:0]\temp_outputs[3] ;   // c:/users/yisong/documents/new/mlp/test.vhd(92[8:20])
    wire [31:0]\hidden_outputs[3] ;   // c:/users/yisong/documents/new/mlp/test.vhd(91[8:22])
    wire [31:0]\temp_outputs[2] ;   // c:/users/yisong/documents/new/mlp/test.vhd(92[8:20])
    wire [31:0]\hidden_outputs[2] ;   // c:/users/yisong/documents/new/mlp/test.vhd(91[8:22])
    wire [31:0]f;   // c:/users/yisong/documents/new/mlp/test.vhd(171[8:9])
    wire [31:0]numL;   // c:/users/yisong/documents/new/mlp/test.vhd(169[8:12])
    wire [31:0]o;   // c:/users/yisong/documents/new/mlp/test.vhd(166[14:15])
    wire mlp_ready;   // c:/users/yisong/documents/new/mlp/main.vhd(303[8:17])
    wire mlp_mode;   // c:/users/yisong/documents/new/mlp/main.vhd(305[8:16])
    wire [31:0]counter;   // c:/users/yisong/documents/new/mlp/test.vhd(167[8:15])
    wire [31:0]i_c;   // c:/users/yisong/documents/new/mlp/test.vhd(166[8:9])
    wire n73801 /* synthesis nomerge= */ ;
    
    wire n23627, n63142, n73806, n62677;
    wire [31:0]n134;
    
    wire n62678, n70697, n24288;
    wire [31:0]n134_adj_403;
    
    wire n62676;
    wire [10:0]n7702;
    
    wire n70712;
    wire [11:0]n13918;
    
    wire n62675, n4593, n62674, n62673, n62672, n62671, n62670;
    wire [31:0]n1027;
    wire [63:0]n2022;
    
    wire n8, n61481;
    wire [10:0]n7729;
    
    wire n5, n62669, n62668, n62667, n62666, n62665, n62664, n73800, 
        n24257;
    wire [31:0]n134_adj_404;
    
    wire n62663, n28, n62662, n62661, n62660, n73807, n23646, 
        n66280, n38, n24, n23647, n63201, n66376, n63210, n73808, 
        n66432, n63239, n66452, n63240, n36, n70731, n4613, n62969, 
        n62659, n62658, n62657, n62656, n62655, n63184, n66340, 
        n62654, n62653, n70848, n3860, n63309, n23658, n62956, 
        n66298, n66454, n62652, n23659, n63188, n62651, n42, n66322, 
        n62650, n62649, n62648, n62647, n66336, n62646, n62645, 
        n66338, n66456, n66334, n63246, n66458, n66460, n66390, 
        n62644, n62643, n66400, n23660, n66300, n66526, n62642, 
        n62641, n62640, n62639, n65, n2239, n62638, n70769, n24023, 
        n62637, n24021, n62636, n70817, n66348, n64, n66474, n62635, 
        n62634, n63058, n62633, n62632, n62631, n23663, n66386, 
        n23664, n63022, n66292, n66468, n23665, n66466, n61484, 
        n12;
    wire [11:0]n3;
    
    wire n61485, n63047, n66530, n66306, n63077, n62613;
    wire [11:0]n54;
    
    wire n62612, n62611, n62610, n60975, n60976, n60974, n62609, 
        n70713, n62608, n62606, n62605, n62604, n62603, n62602, 
        n32, n62600;
    wire [11:0]n3_adj_405;
    wire [11:0]n3_adj_406;
    wire [11:0]n61312;
    
    wire n62599, n62598, n40, n62597, n62596, n70860, n70863, 
        n128, n70857, n70768, n62594;
    wire [11:0]n61292;
    
    wire n62593, n62592, n62591, n62590, n66817, n66247, n65435;
    wire [3:0]n15041;
    
    wire n62589, n61391, n70708, n62588;
    wire [11:0]n61278;
    
    wire n10_adj_71, n4_adj_72, n70809, n46466, n62587, n32_adj_73, 
        n62586, n23234, n44, n62585, n62584, n32_adj_74, n23216, 
        n32_adj_75, n22554, n62583, n31, n34857, n62582, n62581, 
        n66671, n32_adj_76, n23174, n70847;
    wire [31:0]n2448;
    
    wire n1586, n62580, n62579, n22568, n70783, n22745, n62578, 
        n10_adj_77, n62575;
    wire [11:0]n61264;
    
    wire n32_adj_80, n22742, n10_adj_81, n62574, n32_adj_84, n23240, 
        n62573, n17400, n62572, n62571, n40754, n17802, n67260;
    wire [31:0]n1028;
    wire [31:0]n1061;
    
    wire n8_adj_89, n16, n18717, n10_adj_90, n62569;
    wire [11:0]n61250;
    
    wire n62568, n67254, n70842;
    wire [31:0]n3742;
    
    wire n62567, n62566, n62565, n62564, n1585, n70785, n23363, 
        n67252, n67253, n62549;
    wire [11:0]n11102;
    
    wire n32_adj_91, n23237, n62548, n62547, n62546, n62545, n32_adj_92, 
        n23183, n62544, n67541, n67540, n67538, n67537, n67535, 
        n67534, n32_adj_93, n70845, n67532, n23483, n1584, n67531, 
        n67529, n67528, n70786, n23104, n23327, n23330, n1583, 
        n67526, n70861, n1582, n23977, n67525, n67523, n67522, 
        n67520, n67519, n67517, n67516, n32_adj_94, n23297, n81, 
        n23339, n67514, n70787, n22937, n67513, n67511, n32_adj_95, 
        n67510, n67508, n67507, n23186, n67505, n67504, n67502, 
        n67501, n67499, n32_adj_96, n67498, n23321, n67496, n67495, 
        n67493, n32_adj_97, n67492, n67490, n67489, n67487, n22772, 
        n67486, n32_adj_98, n22775, n67484, n67483, n32_adj_99, 
        n70812, n22276, n70736, n23516, n32_adj_100, n23513, n32_adj_101, 
        n22799, n32_adj_102, n23507, n32_adj_103, n23510, n67481, 
        n67480, n67478, n67477, n2664;
    wire [31:0]n134_adj_407;
    
    wire n67475, n67474, n32_adj_105, n67472, n67471, n22548, n67469, 
        n67468, n67466, n67465, n70789, n23360, n32_adj_106, n22802, 
        n32_adj_107, n23207, n67255, n67256, n67257, n61480, n6_adj_108, 
        n66196, n61483, n67258, n67259, n6_adj_109, n70846, n27496, 
        n3756, n77, n60973, n70791, n22748, n66434, n3921, n67264, 
        n67265, n67266, n61486, n61487, n67267, n67268, n67269, 
        n67463, n67462, n67270, n67271, n67272, n67273, n67274, 
        n67275, n67276, n67277, n67278, n32_adj_110, n23504, n23351, 
        n32_adj_111, n67279, n67280, n67281, n66364, n62986, n66366, 
        n63215, n62983, n66436, n63217, n62981, n66362, n66438, 
        n63219, n66440, n62978, n63221, n62976, n66320, n66442, 
        n63227, n63232, n66396, n66342, n66446, n63235, n62972, 
        n66350, n66368, n62990, n63206, n63203, n63213, n63155, 
        n67282, n67283, n67284, n67285, n67286, n67287, n67460, 
        n67459, n67457, n67456, n67454, n67453, n67451, n63119, 
        n67450, n67448, n67447, n67445, n67444, n67288, n67289, 
        n67290, n67442, n67441, n67439, n67438, n67436, n67435, 
        n67433, n67432, n67430, n67429, n67427, n67426, n23975;
    wire [31:0]n134_adj_408;
    
    wire n63158, n63163, n23680, n24020, n63164, n63167, n66556, 
        n2284, n63255, n2277, n2272, n2269, n70701, n2251, n63041, 
        n2242, n63238, n63138, n63135, n63018, n70858, n67291, 
        n67292, n67293, n67294, n67295, n67296, n4923, n62897, 
        n67297, n67298, n67299, n67300, n67301, n67302, n67303, 
        n67304, n67305, n67306, n67307, n67308, n70723, n67309, 
        n67310, n67311, n67312, n67313, n67314, n67315, n67316, 
        n67317, n67318, n67319, n67320, n67321, n67322, n67323, 
        n67324, n67325, n67326, n23968, n67327, n67328, n67329, 
        n67330, n67331, n67332, n67333, n67334, n67335, n67336, 
        n67337, n67338, n67339, n67340, n67341, n67342, n67343, 
        n67344, n67345, n67346, n67347, n67348, n67349, n67350, 
        n63295, n63159, n63254, n70695;
    wire [31:0]n134_adj_409;
    
    wire n67351, n67352, n67353, n67354, n67355, n67356, n67357, 
        n67358, n67359, n67360, n67361, n67362, n67424, n67423, 
        n67421, n67420, n67418, n67417, n67415, n67414, n67412, 
        n67411, n67409, n67408, n67406, n67405, n67363, n67364, 
        n67365, n67366, n67367, n67368, n67369, n67370, n67371, 
        n67403, n67402, n22733, n10_adj_182, n62951, n23282, n67372, 
        n67373, n67374, n67375, n67376, n67377, n67378, n67379, 
        n67380, n10_adj_183, n63065, n23369, n10_adj_185, n66384, 
        n22739, n10_adj_186, n62953, n22913, n10_adj_187, n66408, 
        n22545, n10_adj_188, n66326, n23261, n10_adj_189, n66498, 
        n23447, n10_adj_190, n66360, n67381, n67382, n67383, n23366, 
        n10_adj_191, n63190, n22916, n10_adj_192, n63014, n22928, 
        n10_adj_193, n66318, n23192, n67384, n67385, n67386, n67387, 
        n67388, n67389, n10_adj_194, n66302, n22943, n10_adj_195, 
        n66270, n23354, n10_adj_196, n66388, n23519, n10_adj_199, 
        n66330, n22946, n10_adj_205, n66398, n22940, n10_adj_207, 
        n66276, n22563, n10_adj_222, n66536, n22760, n10_adj_224, 
        n66462, n22551, n10_adj_225, n66268, n22778, n10_adj_226, 
        n66450, n23198, n10_adj_227, n66286, n23138, n10_adj_228, 
        n66424, n22811, n10_adj_229, n66550, n23531, n10_adj_230, 
        n66328, n23318, n10_adj_231, n66546, n22577, n10_adj_232, 
        n62864, n22625, n10_adj_233, n66516, n23492, n10_adj_234, 
        n66344, n22736, n10_adj_235, n66470, n23273, n10_adj_236, 
        n66282, n8_adj_237, n16_adj_238, n17745, n10_adj_239, n67542, 
        n63021, n8_adj_240, n16_adj_241, n17726, n10_adj_242, n67539, 
        n63151;
    wire [31:0]n4478;
    
    wire n70843, n8_adj_243, n67536, n6_adj_244, n36_adj_245, n22931, 
        n10_adj_246, n38_adj_247, n22424, n66484, n8_adj_248, n67530, 
        n6_adj_249, n36_adj_250, n22934, n10_adj_251, n38_adj_252, 
        n66310, n67390, n67391, n67392, n67434, n70859, n8_adj_253, 
        n67527, n6_adj_254, n36_adj_255, n22925, n10_adj_256, n38_adj_257, 
        n66412, n70724, n35, n8_adj_258, n67524, n6_adj_259, n36_adj_260, 
        n22922, n10_adj_261, n38_adj_262, n66404, n32_adj_263, n67393, 
        n67394, n67395, n67518, n22805, n10_adj_264, n16_adj_265, 
        n17644, n12_adj_266, n22919, n63015, n8_adj_267, n16_adj_268, 
        n17638, n10_adj_269, n67515, n63157, n32_adj_270, n8_adj_271, 
        n16_adj_272, n17634, n10_adj_273, n67512, n63161, n8_adj_274, 
        n23501, n16_adj_275, n17619, n10_adj_276, n67509, n63160, 
        n8_adj_277, n16_adj_278, n17405, n10_adj_279, n32_adj_280, 
        n22808, n32_adj_281, n23498, n67506, n63245, n32_adj_282, 
        n22868, n32_adj_283, n23414, n8_adj_284, n67396, n67397, 
        n67398, n32_adj_285, n16_adj_286, n23393, n17365, n10_adj_287, 
        n67503, n32_adj_289, n10_adj_290, n23396, n63165, n8_adj_291, 
        n66528, n66548, n63002, n66420, n66422, n63000, n66428, 
        n66426, n62988, n63207, n66444, n63024, n63027, n66374, 
        n62875, n63223, n63224, n63049, n66356, n62975, n66402, 
        n66448, n63046, n62971, n66346, n66312, n63095, n63052, 
        n66538, n63060, n66284, n62912, n66278, n66514, n63076, 
        n62909, n66540, n66542, n62907, n62855, n66314, n66518, 
        n66562, n62905, n66520, n66410, n66308, n66370, n66382, 
        n63194, n66414, n66380, n66416, n63197, n63004, n66378, 
        n66418, n66332, n62899, n66430, n66324, n66296, n62932, 
        n66492, n63093, n66500, n63094, n62925, n66502, n66304, 
        n63091, n66504, n66272, n62922, n66274, n63192, n66506, 
        n63083, n62920, n66290, n66406, n63078, n66508, n66294, 
        n62916, n63085, n66510, n66288, n66266, n62914, n63080, 
        n66512, n16_adj_292, n17345, n10_adj_293, n67500, n63253, 
        n8_adj_294, n67399, n67400, n67401, n16_adj_295, n17309, 
        n10_adj_296, n67497, n63153, n8_adj_297, n16_adj_298, n17887, 
        n10_adj_299, n67494, n63146, n8_adj_300, n66472, n66486, 
        n62949, n62948, n66476, n63168, n62946, n66394, n66552, 
        n66478, n66392, n62944, n63173, n66554, n66480, n63199, 
        n62942, n66372, n66482, n66496, n62940, n66358, n62938, 
        n66354, n62937, n66352, n66488, n66544, n62934, n63252, 
        n66490, n63118, n63117, n63132, n63134, n63149, n63256, 
        n63137, n63136, n63143, n63140, n63141, n63144, n63196, 
        n63145, n23357, n67404, n16_adj_301, n17567, n10_adj_302, 
        n67491, n67407, n8_adj_303, n16_adj_304, n17891, n10_adj_305, 
        n67488, n67410, n70725, n8_adj_306, n16_adj_307, n17895, 
        n10_adj_308, n67485, n22607, n22610, n67413, n67416, n8_adj_309, 
        n16_adj_310, n67419, n67422, n17899, n10_adj_311, n67482, 
        n39, n51, n46, n8_adj_312, n56_adj_313, n16_adj_314, n17901, 
        n10_adj_315, n67479, n42_adj_316, n1, n60_adj_317;
    wire [11:0]n13947;
    
    wire n41, n8_adj_318, n50, n58_adj_319, n62_adj_320, n49, n16_adj_321, 
        n17905, n10_adj_322, n67476, n8_adj_323, n67425, n16_adj_324, 
        n17909, n10_adj_325, n67473, n8_adj_326, n16_adj_327, n17911, 
        n10_adj_328, n67470, n67443, n8_adj_330, n23525, n16_adj_331, 
        n17881, n10_adj_332, n67467, n23528, n8_adj_333, n16_adj_334, 
        n17919, n10_adj_335, n67464, n8_adj_336, n16_adj_337, n17921, 
        n10_adj_338, n67461, n8_adj_339, n16_adj_340, n17925, n10_adj_341, 
        n67458, n8_adj_342, n16_adj_343, n18121, n10_adj_344, n67455, 
        n67440, n8_adj_345, n23, n1423, n16_adj_346, n18119, n10_adj_347, 
        n67452, n70700, n23345, n23348, n22682, n23189, n22685, 
        n23534, n3922, n22688, n67428, n23495, n22691, n23465, 
        n22694, n23459, n22697, n23417, n22700, n67431, n23405, 
        n67437, n22703, n23390, n67446, n67449, n22706, n23315, 
        n23312, n22712, n23309, n22715, n23306, n23303, n22718, 
        n23300, n22721, n22724, n22727, n23291, n22730, n22637, 
        n23270, n22640, n23267, n23264, n22643, n23258, n22646, 
        n23255, n22649, n23252, n22652, n23246, n22655, n23243, 
        n22658, n23372, n23231, n22661, n23228, n22664, n23225, 
        n23222, n22667, n22670, n23210, n22673, n23201, n22676, 
        n22679, n23195, n60990, n22598, n22874, n22601, n22841, 
        n22898, n23387, n22901, n23384, n22904, n23381, n22907, 
        n23378, n23375, n23420, n22826, n22910, n22613, n22616, 
        n67521, n22709, n22619, n22583, n22569, n22622, n22557, 
        n23294, n22628, n23288, n22631, n23279, n22634, n23276, 
        n23249, n22560, n23219, n23213, n23177, n23489, n22814, 
        n23171, n67533, n22820, n23168, n22829, n23462, n23180, 
        n23456, n23453, n22589, n23399, n23135, n23132, n22592, 
        n60989, n23411, n22871, n22883, n22880, n22889, n22886, 
        n22892, n22895, n23129, n22595, n70864, n8_adj_349, n38_adj_350, 
        n17650, n10_adj_351, n8_adj_352, n38_adj_353, n17704, n10_adj_354, 
        n60988, n60987, n22865, n60986, n6_adj_355, n7_adj_356, 
        n6_adj_357, n7_adj_358, n6_adj_359, n7_adj_360, n6_adj_361, 
        n7_adj_362, n38_adj_363, n52, n46_adj_364, n56_adj_365, n42_adj_366, 
        n54_adj_367, n60_adj_368, n41_adj_369, n50_adj_370, n58_adj_371, 
        n62_adj_372, n49_adj_373, n60985, n6_adj_374, n7_adj_375, 
        n66837, n66975, n66845, n66979, n67013, n66847, n66987, 
        n66983, n66985, n67029, n67019, n67037, n63590, n6_adj_376, 
        n7_adj_377, n6_adj_378, n7_adj_379, n12_adj_380, n6_adj_381, 
        n7_adj_382, n6_adj_383, n7_adj_384, n40_adj_385, n50_adj_386, 
        n36_adj_387, n48, n32_adj_388, n46_adj_389, n44_adj_390, n52_adj_391, 
        n54_adj_392, n53, n55_adj_393, n60984, n62189, n62188, n62187, 
        n62186, n62185, n62184, n62183, n62182, n62181, n62180, 
        n22793, n22796, n62179, n62178, n62177, n22784, n22787, 
        n23123, n23126, n23114, n23117, n62176, n62175, n23105, 
        n23108, n62174, n60983, n23096, n23099, n23087, n23090, 
        n23078, n23081, n23069, n23072, n23060, n23063, n23051, 
        n23054, n60982, n23033, n23036, n23042, n23045, n23024, 
        n23027, n23006, n23009, n23015, n23018, n22997, n23000, 
        n22988, n22991, n22979, n22982, n60981, n22766, n22769, 
        n22970, n22973, n22961, n22964, n70813, n6_adj_394, n4_adj_395, 
        n4_adj_396, n22754, n22757;
    wire [31:0]n3998;
    
    wire n22952, n22955, n60980, n6_adj_397, n7_adj_398, n6_adj_399, 
        n7_adj_400, n23426, n23402, n23408, n22877, n23423, n23480, 
        n22817, n23486, n22823, n23471, n22586, n23477, n23468, 
        n60979, n22835, n23474, n70862, n22832, n23450, n22838, 
        n22844, n23444, n22847, n23441, n22850, n23438, n22853, 
        n22856, n23432, n23429, n22862, n23435, n61477, n67623, 
        n22859, n6_adj_401, n61478, n2, n60978, n61479, n8_adj_402, 
        n62765, n62764, n62763, n62762, n62761, n62760, n61482, 
        n60977, n63026, n62711, n62710, n62709, n66887, n62708, 
        n62707, n62706, n62705, n62704, n62703, n62702, n62701, 
        n62700, n62699, n62698, n62697, n62696, n62694, n62693, 
        n62692, n62691, n62690, n62689, n62688, n62687, n62686, 
        n62685, n62684, n62683, n62682, n62681, n62680;
    
    FD1P3AX sram_addr_i0_i0 (.D(n63142), .SP(n23627), .CK(clock), .Q(sram_address_B[0]));
    defparam sram_addr_i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i23 (.D(\hidden_outputs[1] [23]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [23]));
    defparam temp_outputs_1__i0_i23.GSR = "DISABLED";
    CCU2D h_4657_add_4_31 (.A0(h[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62677), 
          .COUT(n62678), .S0(n134[29]), .S1(n134[30]));
    defparam h_4657_add_4_31.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_31.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_31.INJECT1_0 = "NO";
    defparam h_4657_add_4_31.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i22 (.D(\hidden_outputs[1] [22]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [22]));
    defparam temp_outputs_1__i0_i22.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i21 (.D(\hidden_outputs[1] [21]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [21]));
    defparam temp_outputs_1__i0_i21.GSR = "DISABLED";
    FD1P3IX n_4659__i16 (.D(n134_adj_403[16]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[16]));
    defparam n_4659__i16.GSR = "DISABLED";
    CCU2D h_4657_add_4_29 (.A0(h[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62676), 
          .COUT(n62677), .S0(n134[27]), .S1(n134[28]));
    defparam h_4657_add_4_29.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_29.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_29.INJECT1_0 = "NO";
    defparam h_4657_add_4_29.INJECT1_1 = "NO";
    LUT4 mux_4578_i5_3_lut (.A(n7702[3]), .B(h[4]), .C(n70712), .Z(n13918[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4578_i5_3_lut.init = 16'hcaca;
    FD1P3IX n_4659__i15 (.D(n134_adj_403[15]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[15]));
    defparam n_4659__i15.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i5 (.D(\hidden_outputs[0] [5]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [5]));
    defparam temp_outputs_0__i0_i5.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i16 (.D(\hidden_outputs[0] [16]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [16]));
    defparam temp_outputs_0__i0_i16.GSR = "DISABLED";
    CCU2D h_4657_add_4_27 (.A0(h[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62675), 
          .COUT(n62676), .S0(n134[25]), .S1(n134[26]));
    defparam h_4657_add_4_27.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_27.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_27.INJECT1_0 = "NO";
    defparam h_4657_add_4_27.INJECT1_1 = "NO";
    FD1P3IX n_4659__i14 (.D(n134_adj_403[14]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[14]));
    defparam n_4659__i14.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i25 (.D(\hidden_outputs[1] [25]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [25]));
    defparam temp_outputs_1__i0_i25.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i15 (.D(\hidden_outputs[0] [15]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [15]));
    defparam temp_outputs_0__i0_i15.GSR = "DISABLED";
    FD1P3IX n_4659__i13 (.D(n134_adj_403[13]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[13]));
    defparam n_4659__i13.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i4 (.D(\hidden_outputs[0] [4]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [4]));
    defparam temp_outputs_0__i0_i4.GSR = "DISABLED";
    FD1P3AX weight_i0_i0 (.D(sram_output_B[0]), .SP(n4593), .CK(clock), 
            .Q(weight[0]));
    defparam weight_i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i20 (.D(\hidden_outputs[1] [20]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [20]));
    defparam temp_outputs_1__i0_i20.GSR = "DISABLED";
    CCU2D h_4657_add_4_25 (.A0(h[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62674), 
          .COUT(n62675), .S0(n134[23]), .S1(n134[24]));
    defparam h_4657_add_4_25.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_25.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_25.INJECT1_0 = "NO";
    defparam h_4657_add_4_25.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_23 (.A0(h[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62673), 
          .COUT(n62674), .S0(n134[21]), .S1(n134[22]));
    defparam h_4657_add_4_23.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_23.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_23.INJECT1_0 = "NO";
    defparam h_4657_add_4_23.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i19 (.D(\hidden_outputs[1] [19]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [19]));
    defparam temp_outputs_1__i0_i19.GSR = "DISABLED";
    CCU2D h_4657_add_4_21 (.A0(h[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62672), 
          .COUT(n62673), .S0(n134[19]), .S1(n134[20]));
    defparam h_4657_add_4_21.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_21.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_21.INJECT1_0 = "NO";
    defparam h_4657_add_4_21.INJECT1_1 = "NO";
    FD1P3AX e_i0_i0 (.D(float_alu_c[0]), .SP(n4599), .CK(clock), .Q(e[0]));
    defparam e_i0_i0.GSR = "DISABLED";
    CCU2D h_4657_add_4_19 (.A0(h[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62671), 
          .COUT(n62672), .S0(n134[17]), .S1(n134[18]));
    defparam h_4657_add_4_19.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_19.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_19.INJECT1_0 = "NO";
    defparam h_4657_add_4_19.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_17 (.A0(h[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62670), 
          .COUT(n62671), .S0(n134[15]), .S1(n134[16]));
    defparam h_4657_add_4_17.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_17.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_17.INJECT1_0 = "NO";
    defparam h_4657_add_4_17.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i18 (.D(\hidden_outputs[1] [18]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [18]));
    defparam temp_outputs_1__i0_i18.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i17 (.D(\hidden_outputs[1] [17]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [17]));
    defparam temp_outputs_1__i0_i17.GSR = "DISABLED";
    DPR16X4C inputs1 (.DI0(sram_output_B[24]), .DI1(sram_output_B[25]), 
            .DI2(sram_output_B[26]), .DI3(sram_output_B[27]), .WAD0(addr[0]), 
            .WAD1(addr[1]), .WAD2(addr[2]), .WAD3(GND_net), .WCK(clock), 
            .WRE(n15113), .RAD0(i[0]), .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), 
            .DO0(n1027[24]), .DO1(n1027[25]), .DO2(n1027[26]), .DO3(n1027[27]));
    defparam inputs1.initval = "0x0000000000000000";
    FD1P3AX temp_outputs_1__i0_i16 (.D(\hidden_outputs[1] [16]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [16]));
    defparam temp_outputs_1__i0_i16.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i15 (.D(\hidden_outputs[1] [15]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [15]));
    defparam temp_outputs_1__i0_i15.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i14 (.D(\hidden_outputs[1] [14]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [14]));
    defparam temp_outputs_1__i0_i14.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i13 (.D(\hidden_outputs[1] [13]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [13]));
    defparam temp_outputs_1__i0_i13.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i0 (.D(\hidden_outputs[4] [0]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[4] [0]));
    defparam temp_outputs_4__i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i12 (.D(\hidden_outputs[1] [12]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [12]));
    defparam temp_outputs_1__i0_i12.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i11 (.D(\hidden_outputs[1] [11]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [11]));
    defparam temp_outputs_1__i0_i11.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i0 (.D(\hidden_outputs[3] [0]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[3] [0]));
    defparam temp_outputs_3__i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i0 (.D(\hidden_outputs[2] [0]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [0]));
    defparam temp_outputs_2__i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i0 (.D(\hidden_outputs[1] [0]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [0]));
    defparam temp_outputs_1__i0_i0.GSR = "DISABLED";
    LUT4 i3_3_lut (.A(n2022[10]), .B(n2022[7]), .C(n2022[32]), .Z(n8)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i3_3_lut.init = 16'hfefe;
    FD1P3AX temp_outputs_0__i0_i0 (.D(\hidden_outputs[0] [0]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [0]));
    defparam temp_outputs_0__i0_i0.GSR = "DISABLED";
    FD1P3AX f_i0_i0 (.D(float_alu_c[0]), .SP(n4617), .CK(clock), .Q(f[0]));
    defparam f_i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i10 (.D(\hidden_outputs[1] [10]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [10]));
    defparam temp_outputs_1__i0_i10.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i3 (.D(\hidden_outputs[0] [3]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [3]));
    defparam temp_outputs_0__i0_i3.GSR = "DISABLED";
    FD1P3IX n_4659__i12 (.D(n134_adj_403[12]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[12]));
    defparam n_4659__i12.GSR = "DISABLED";
    FD1P3IX n_4659__i11 (.D(n134_adj_403[11]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[11]));
    defparam n_4659__i11.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i9 (.D(\hidden_outputs[1] [9]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [9]));
    defparam temp_outputs_1__i0_i9.GSR = "DISABLED";
    CCU2D add_4597_12 (.A0(i[10]), .B0(h[11]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n61481), 
          .S0(n7729[10]));
    defparam add_4597_12.INIT0 = 16'h5666;
    defparam add_4597_12.INIT1 = 16'h0000;
    defparam add_4597_12.INJECT1_0 = "NO";
    defparam add_4597_12.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(numL[0]), .B(n14054), .Z(n5)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX n_4659__i10 (.D(n134_adj_403[10]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[10]));
    defparam n_4659__i10.GSR = "DISABLED";
    FD1P3IX n_4659__i9 (.D(n134_adj_403[9]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[9]));
    defparam n_4659__i9.GSR = "DISABLED";
    FD1P3IX n_4659__i8 (.D(n134_adj_403[8]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[8]));
    defparam n_4659__i8.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i8 (.D(\hidden_outputs[1] [8]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [8]));
    defparam temp_outputs_1__i0_i8.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i7 (.D(\hidden_outputs[1] [7]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [7]));
    defparam temp_outputs_1__i0_i7.GSR = "DISABLED";
    FD1P3IX n_4659__i7 (.D(n134_adj_403[7]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[7]));
    defparam n_4659__i7.GSR = "DISABLED";
    FD1P3IX n_4659__i6 (.D(n134_adj_403[6]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[6]));
    defparam n_4659__i6.GSR = "DISABLED";
    FD1P3IX n_4659__i5 (.D(n134_adj_403[5]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[5]));
    defparam n_4659__i5.GSR = "DISABLED";
    LUT4 i27931_4_lut (.A(n2022[29]), .B(n70822), .C(n8), .D(n2022[1]), 
         .Z(n23627)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i27931_4_lut.init = 16'hccc8;
    CCU2D h_4657_add_4_15 (.A0(h[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62669), 
          .COUT(n62670), .S0(n134[13]), .S1(n134[14]));
    defparam h_4657_add_4_15.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_15.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_15.INJECT1_0 = "NO";
    defparam h_4657_add_4_15.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_13 (.A0(h[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62668), 
          .COUT(n62669), .S0(n134[11]), .S1(n134[12]));
    defparam h_4657_add_4_13.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_13.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_13.INJECT1_0 = "NO";
    defparam h_4657_add_4_13.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_11 (.A0(h[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62667), 
          .COUT(n62668), .S0(n134[9]), .S1(n134[10]));
    defparam h_4657_add_4_11.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_11.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_11.INJECT1_0 = "NO";
    defparam h_4657_add_4_11.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_9 (.A0(h[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62666), 
          .COUT(n62667), .S0(n134[7]), .S1(n134[8]));
    defparam h_4657_add_4_9.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_9.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_9.INJECT1_0 = "NO";
    defparam h_4657_add_4_9.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_7 (.A0(h[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62665), 
          .COUT(n62666), .S0(n134[5]), .S1(n134[6]));
    defparam h_4657_add_4_7.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_7.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_7.INJECT1_0 = "NO";
    defparam h_4657_add_4_7.INJECT1_1 = "NO";
    FD1P3IX n_4659__i4 (.D(n134_adj_403[4]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[4]));
    defparam n_4659__i4.GSR = "DISABLED";
    FD1P3IX n_4659__i3 (.D(n134_adj_403[3]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[3]));
    defparam n_4659__i3.GSR = "DISABLED";
    CCU2D h_4657_add_4_5 (.A0(h[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62664), 
          .COUT(n62665), .S0(n134[3]), .S1(n134[4]));
    defparam h_4657_add_4_5.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_5.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_5.INJECT1_0 = "NO";
    defparam h_4657_add_4_5.INJECT1_1 = "NO";
    FD1P3IX n_4659__i2 (.D(n134_adj_403[2]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[2]));
    defparam n_4659__i2.GSR = "DISABLED";
    FD1P3IX n_4659__i17 (.D(n134_adj_403[17]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[17]));
    defparam n_4659__i17.GSR = "DISABLED";
    FD1P3IX n_4659__i1 (.D(n134_adj_403[1]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[1]));
    defparam n_4659__i1.GSR = "DISABLED";
    FD1P3IX o_4661__i31 (.D(n134_adj_404[31]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[31]));
    defparam o_4661__i31.GSR = "DISABLED";
    CCU2D h_4657_add_4_3 (.A0(h[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62663), 
          .COUT(n62664), .S0(n134[1]), .S1(n134[2]));
    defparam h_4657_add_4_3.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_3.INIT1 = 16'hfaaa;
    defparam h_4657_add_4_3.INJECT1_0 = "NO";
    defparam h_4657_add_4_3.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_0__i0_i14 (.D(\hidden_outputs[0] [14]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[0] [14]));
    defparam temp_outputs_0__i0_i14.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i6 (.D(\hidden_outputs[1] [6]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [6]));
    defparam temp_outputs_1__i0_i6.GSR = "DISABLED";
    CCU2D h_4657_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62663), 
          .S1(n134[0]));
    defparam h_4657_add_4_1.INIT0 = 16'hF000;
    defparam h_4657_add_4_1.INIT1 = 16'h0555;
    defparam h_4657_add_4_1.INJECT1_0 = "NO";
    defparam h_4657_add_4_1.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i5 (.D(\hidden_outputs[1] [5]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [5]));
    defparam temp_outputs_1__i0_i5.GSR = "DISABLED";
    LUT4 i5_2_lut (.A(numL[10]), .B(numL[17]), .Z(n28)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    FD1P3AX temp_outputs_1__i0_i4 (.D(\hidden_outputs[1] [4]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [4]));
    defparam temp_outputs_1__i0_i4.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i3 (.D(\hidden_outputs[1] [3]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [3]));
    defparam temp_outputs_1__i0_i3.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i2 (.D(\hidden_outputs[1] [2]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [2]));
    defparam temp_outputs_1__i0_i2.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i1 (.D(\hidden_outputs[1] [1]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[1] [1]));
    defparam temp_outputs_1__i0_i1.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i31 (.D(\hidden_outputs[2] [31]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [31]));
    defparam temp_outputs_2__i0_i31.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i30 (.D(\hidden_outputs[2] [30]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [30]));
    defparam temp_outputs_2__i0_i30.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i29 (.D(\hidden_outputs[2] [29]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [29]));
    defparam temp_outputs_2__i0_i29.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i28 (.D(\hidden_outputs[2] [28]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [28]));
    defparam temp_outputs_2__i0_i28.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i27 (.D(\hidden_outputs[2] [27]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [27]));
    defparam temp_outputs_2__i0_i27.GSR = "DISABLED";
    CCU2D n_4659_add_4_33 (.A0(n[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62662), 
          .S0(n134_adj_403[31]));
    defparam n_4659_add_4_33.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_33.INIT1 = 16'h0000;
    defparam n_4659_add_4_33.INJECT1_0 = "NO";
    defparam n_4659_add_4_33.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_2__i0_i26 (.D(\hidden_outputs[2] [26]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [26]));
    defparam temp_outputs_2__i0_i26.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i25 (.D(\hidden_outputs[2] [25]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [25]));
    defparam temp_outputs_2__i0_i25.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i24 (.D(\hidden_outputs[2] [24]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [24]));
    defparam temp_outputs_2__i0_i24.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i23 (.D(\hidden_outputs[2] [23]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [23]));
    defparam temp_outputs_2__i0_i23.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i22 (.D(\hidden_outputs[2] [22]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [22]));
    defparam temp_outputs_2__i0_i22.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i21 (.D(\hidden_outputs[2] [21]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [21]));
    defparam temp_outputs_2__i0_i21.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i20 (.D(\hidden_outputs[2] [20]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [20]));
    defparam temp_outputs_2__i0_i20.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i19 (.D(\hidden_outputs[2] [19]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [19]));
    defparam temp_outputs_2__i0_i19.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i18 (.D(\hidden_outputs[2] [18]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [18]));
    defparam temp_outputs_2__i0_i18.GSR = "DISABLED";
    CCU2D n_4659_add_4_31 (.A0(n[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62661), 
          .COUT(n62662), .S0(n134_adj_403[29]), .S1(n134_adj_403[30]));
    defparam n_4659_add_4_31.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_31.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_31.INJECT1_0 = "NO";
    defparam n_4659_add_4_31.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_29 (.A0(n[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62660), 
          .COUT(n62661), .S0(n134_adj_403[27]), .S1(n134_adj_403[28]));
    defparam n_4659_add_4_29.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_29.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_29.INJECT1_0 = "NO";
    defparam n_4659_add_4_29.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_2__i0_i17 (.D(\hidden_outputs[2] [17]), .SP(n73806), 
            .CK(clock), .Q(\temp_outputs[2] [17]));
    defparam temp_outputs_2__i0_i17.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i16 (.D(\hidden_outputs[2] [16]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [16]));
    defparam temp_outputs_2__i0_i16.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i15 (.D(\hidden_outputs[2] [15]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [15]));
    defparam temp_outputs_2__i0_i15.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i14 (.D(\hidden_outputs[2] [14]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [14]));
    defparam temp_outputs_2__i0_i14.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i13 (.D(\hidden_outputs[2] [13]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [13]));
    defparam temp_outputs_2__i0_i13.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i12 (.D(\hidden_outputs[2] [12]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [12]));
    defparam temp_outputs_2__i0_i12.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i11 (.D(\hidden_outputs[2] [11]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [11]));
    defparam temp_outputs_2__i0_i11.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i10 (.D(\hidden_outputs[2] [10]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [10]));
    defparam temp_outputs_2__i0_i10.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i9 (.D(\hidden_outputs[2] [9]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [9]));
    defparam temp_outputs_2__i0_i9.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i8 (.D(\hidden_outputs[2] [8]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [8]));
    defparam temp_outputs_2__i0_i8.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i7 (.D(\hidden_outputs[2] [7]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [7]));
    defparam temp_outputs_2__i0_i7.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i6 (.D(\hidden_outputs[2] [6]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [6]));
    defparam temp_outputs_2__i0_i6.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i5 (.D(\hidden_outputs[2] [5]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [5]));
    defparam temp_outputs_2__i0_i5.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i4 (.D(\hidden_outputs[2] [4]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [4]));
    defparam temp_outputs_2__i0_i4.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i3 (.D(\hidden_outputs[2] [3]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [3]));
    defparam temp_outputs_2__i0_i3.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i2 (.D(\hidden_outputs[2] [2]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [2]));
    defparam temp_outputs_2__i0_i2.GSR = "DISABLED";
    FD1P3AX temp_outputs_2__i0_i1 (.D(\hidden_outputs[2] [1]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[2] [1]));
    defparam temp_outputs_2__i0_i1.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i31 (.D(\hidden_outputs[3] [31]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [31]));
    defparam temp_outputs_3__i0_i31.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i30 (.D(\hidden_outputs[3] [30]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [30]));
    defparam temp_outputs_3__i0_i30.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i29 (.D(\hidden_outputs[3] [29]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [29]));
    defparam temp_outputs_3__i0_i29.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i28 (.D(\hidden_outputs[3] [28]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [28]));
    defparam temp_outputs_3__i0_i28.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i27 (.D(\hidden_outputs[3] [27]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [27]));
    defparam temp_outputs_3__i0_i27.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i0 (.D(n66280), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [0]));
    defparam output_outputs_0__i0_i0.GSR = "DISABLED";
    LUT4 i15_4_lut (.A(numL[28]), .B(numL[2]), .C(numL[5]), .D(numL[11]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_1 (.A(numL[30]), .B(numL[15]), .Z(n24)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_1.init = 16'heeee;
    FD1P3AX temp_outputs_3__i0_i26 (.D(\hidden_outputs[3] [26]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [26]));
    defparam temp_outputs_3__i0_i26.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i25 (.D(\hidden_outputs[3] [25]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [25]));
    defparam temp_outputs_3__i0_i25.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i24 (.D(\hidden_outputs[3] [24]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [24]));
    defparam temp_outputs_3__i0_i24.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i23 (.D(\hidden_outputs[3] [23]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [23]));
    defparam temp_outputs_3__i0_i23.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i22 (.D(\hidden_outputs[3] [22]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [22]));
    defparam temp_outputs_3__i0_i22.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i21 (.D(\hidden_outputs[3] [21]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [21]));
    defparam temp_outputs_3__i0_i21.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i20 (.D(\hidden_outputs[3] [20]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [20]));
    defparam temp_outputs_3__i0_i20.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i19 (.D(\hidden_outputs[3] [19]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [19]));
    defparam temp_outputs_3__i0_i19.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i18 (.D(\hidden_outputs[3] [18]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [18]));
    defparam temp_outputs_3__i0_i18.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i17 (.D(\hidden_outputs[3] [17]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [17]));
    defparam temp_outputs_3__i0_i17.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i16 (.D(\hidden_outputs[3] [16]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [16]));
    defparam temp_outputs_3__i0_i16.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i15 (.D(\hidden_outputs[3] [15]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [15]));
    defparam temp_outputs_3__i0_i15.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i14 (.D(\hidden_outputs[3] [14]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [14]));
    defparam temp_outputs_3__i0_i14.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i13 (.D(\hidden_outputs[3] [13]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [13]));
    defparam temp_outputs_3__i0_i13.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i12 (.D(\hidden_outputs[3] [12]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [12]));
    defparam temp_outputs_3__i0_i12.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i11 (.D(\hidden_outputs[3] [11]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [11]));
    defparam temp_outputs_3__i0_i11.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i10 (.D(\hidden_outputs[3] [10]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [10]));
    defparam temp_outputs_3__i0_i10.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i9 (.D(\hidden_outputs[3] [9]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [9]));
    defparam temp_outputs_3__i0_i9.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i8 (.D(\hidden_outputs[3] [8]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [8]));
    defparam temp_outputs_3__i0_i8.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i7 (.D(\hidden_outputs[3] [7]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [7]));
    defparam temp_outputs_3__i0_i7.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i6 (.D(\hidden_outputs[3] [6]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [6]));
    defparam temp_outputs_3__i0_i6.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i5 (.D(\hidden_outputs[3] [5]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [5]));
    defparam temp_outputs_3__i0_i5.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i4 (.D(\hidden_outputs[3] [4]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [4]));
    defparam temp_outputs_3__i0_i4.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i3 (.D(\hidden_outputs[3] [3]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [3]));
    defparam temp_outputs_3__i0_i3.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i31 (.D(n63201), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [31]));
    defparam output_outputs_1__i0_i31.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i2 (.D(\hidden_outputs[3] [2]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [2]));
    defparam temp_outputs_3__i0_i2.GSR = "DISABLED";
    FD1P3AX temp_outputs_3__i0_i1 (.D(\hidden_outputs[3] [1]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[3] [1]));
    defparam temp_outputs_3__i0_i1.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i30 (.D(n66376), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [30]));
    defparam output_outputs_1__i0_i30.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i31 (.D(\hidden_outputs[4] [31]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[4] [31]));
    defparam temp_outputs_4__i0_i31.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i30 (.D(\hidden_outputs[4] [30]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[4] [30]));
    defparam temp_outputs_4__i0_i30.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i29 (.D(n63210), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [29]));
    defparam output_outputs_1__i0_i29.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i29 (.D(\hidden_outputs[4] [29]), .SP(n73807), 
            .CK(clock), .Q(\temp_outputs[4] [29]));
    defparam temp_outputs_4__i0_i29.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i28 (.D(\hidden_outputs[4] [28]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [28]));
    defparam temp_outputs_4__i0_i28.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i28 (.D(n66432), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [28]));
    defparam output_outputs_1__i0_i28.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i27 (.D(\hidden_outputs[4] [27]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [27]));
    defparam temp_outputs_4__i0_i27.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i26 (.D(\hidden_outputs[4] [26]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [26]));
    defparam temp_outputs_4__i0_i26.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i25 (.D(\hidden_outputs[4] [25]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [25]));
    defparam temp_outputs_4__i0_i25.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i24 (.D(\hidden_outputs[4] [24]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [24]));
    defparam temp_outputs_4__i0_i24.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i23 (.D(\hidden_outputs[4] [23]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [23]));
    defparam temp_outputs_4__i0_i23.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i22 (.D(\hidden_outputs[4] [22]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [22]));
    defparam temp_outputs_4__i0_i22.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i27 (.D(n63239), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [27]));
    defparam output_outputs_1__i0_i27.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i26 (.D(n66452), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [26]));
    defparam output_outputs_1__i0_i26.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i25 (.D(n63240), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [25]));
    defparam output_outputs_1__i0_i25.GSR = "DISABLED";
    LUT4 i13_4_lut (.A(numL[19]), .B(numL[23]), .C(numL[12]), .D(numL[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_rep_910 (.A(n70731), .B(n14054), .C(n4613), 
         .D(numL[31]), .Z(n73808)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_rep_910.init = 16'hf010;
    FD1P3AX output_outputs_1__i0_i24 (.D(n62969), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [24]));
    defparam output_outputs_1__i0_i24.GSR = "DISABLED";
    CCU2D n_4659_add_4_27 (.A0(n[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62659), 
          .COUT(n62660), .S0(n134_adj_403[25]), .S1(n134_adj_403[26]));
    defparam n_4659_add_4_27.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_27.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_27.INJECT1_0 = "NO";
    defparam n_4659_add_4_27.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_25 (.A0(n[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62658), 
          .COUT(n62659), .S0(n134_adj_403[23]), .S1(n134_adj_403[24]));
    defparam n_4659_add_4_25.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_25.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_25.INJECT1_0 = "NO";
    defparam n_4659_add_4_25.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_23 (.A0(n[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62657), 
          .COUT(n62658), .S0(n134_adj_403[21]), .S1(n134_adj_403[22]));
    defparam n_4659_add_4_23.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_23.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_23.INJECT1_0 = "NO";
    defparam n_4659_add_4_23.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_21 (.A0(n[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62656), 
          .COUT(n62657), .S0(n134_adj_403[19]), .S1(n134_adj_403[20]));
    defparam n_4659_add_4_21.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_21.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_21.INJECT1_0 = "NO";
    defparam n_4659_add_4_21.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_4__i0_i21 (.D(\hidden_outputs[4] [21]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [21]));
    defparam temp_outputs_4__i0_i21.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i20 (.D(\hidden_outputs[4] [20]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [20]));
    defparam temp_outputs_4__i0_i20.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i19 (.D(\hidden_outputs[4] [19]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [19]));
    defparam temp_outputs_4__i0_i19.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i18 (.D(\hidden_outputs[4] [18]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [18]));
    defparam temp_outputs_4__i0_i18.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i17 (.D(\hidden_outputs[4] [17]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [17]));
    defparam temp_outputs_4__i0_i17.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i16 (.D(\hidden_outputs[4] [16]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [16]));
    defparam temp_outputs_4__i0_i16.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i15 (.D(\hidden_outputs[4] [15]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [15]));
    defparam temp_outputs_4__i0_i15.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i14 (.D(\hidden_outputs[4] [14]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [14]));
    defparam temp_outputs_4__i0_i14.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i13 (.D(\hidden_outputs[4] [13]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [13]));
    defparam temp_outputs_4__i0_i13.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i12 (.D(\hidden_outputs[4] [12]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [12]));
    defparam temp_outputs_4__i0_i12.GSR = "DISABLED";
    CCU2D n_4659_add_4_19 (.A0(n[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62655), 
          .COUT(n62656), .S0(n134_adj_403[17]), .S1(n134_adj_403[18]));
    defparam n_4659_add_4_19.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_19.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_19.INJECT1_0 = "NO";
    defparam n_4659_add_4_19.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_4__i0_i11 (.D(\hidden_outputs[4] [11]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [11]));
    defparam temp_outputs_4__i0_i11.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i10 (.D(\hidden_outputs[4] [10]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [10]));
    defparam temp_outputs_4__i0_i10.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i9 (.D(\hidden_outputs[4] [9]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [9]));
    defparam temp_outputs_4__i0_i9.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i8 (.D(\hidden_outputs[4] [8]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [8]));
    defparam temp_outputs_4__i0_i8.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i7 (.D(\hidden_outputs[4] [7]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [7]));
    defparam temp_outputs_4__i0_i7.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i6 (.D(\hidden_outputs[4] [6]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [6]));
    defparam temp_outputs_4__i0_i6.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i5 (.D(\hidden_outputs[4] [5]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [5]));
    defparam temp_outputs_4__i0_i5.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i4 (.D(\hidden_outputs[4] [4]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [4]));
    defparam temp_outputs_4__i0_i4.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i3 (.D(\hidden_outputs[4] [3]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [3]));
    defparam temp_outputs_4__i0_i3.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i2 (.D(\hidden_outputs[4] [2]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [2]));
    defparam temp_outputs_4__i0_i2.GSR = "DISABLED";
    FD1P3AX temp_outputs_4__i0_i1 (.D(\hidden_outputs[4] [1]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[4] [1]));
    defparam temp_outputs_4__i0_i1.GSR = "DISABLED";
    FD1P3AX e_i0_i31 (.D(float_alu_c[31]), .SP(n4599), .CK(clock), .Q(e[31]));
    defparam e_i0_i31.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i0 (.D(n63184), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [0]));
    defparam output_outputs_1__i0_i0.GSR = "DISABLED";
    FD1P3AX e_i0_i30 (.D(float_alu_c[30]), .SP(n4599), .CK(clock), .Q(e[30]));
    defparam e_i0_i30.GSR = "DISABLED";
    FD1P3IX o_4661__i30 (.D(n134_adj_404[30]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[30]));
    defparam o_4661__i30.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i23 (.D(n66340), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [23]));
    defparam output_outputs_1__i0_i23.GSR = "DISABLED";
    CCU2D n_4659_add_4_17 (.A0(n[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62654), 
          .COUT(n62655), .S0(n134_adj_403[15]), .S1(n134_adj_403[16]));
    defparam n_4659_add_4_17.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_17.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_17.INJECT1_0 = "NO";
    defparam n_4659_add_4_17.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_15 (.A0(n[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62653), 
          .COUT(n62654), .S0(n134_adj_403[13]), .S1(n134_adj_403[14]));
    defparam n_4659_add_4_15.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_15.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_15.INJECT1_0 = "NO";
    defparam n_4659_add_4_15.INJECT1_1 = "NO";
    FD1P3DX ready_437 (.D(n70848), .SP(n23653), .CK(clock), .CD(SDA_c), 
            .Q(mlp_ready));
    defparam ready_437.GSR = "DISABLED";
    FD1P3DX sram_ready_441 (.D(n3860), .SP(n23655), .CK(clock), .CD(SDA_c), 
            .Q(sram_ready_B));
    defparam sram_ready_441.GSR = "DISABLED";
    FD1S3DX mlp_mode_20 (.D(n63309), .CK(clock), .CD(SDA_c), .Q(mlp_mode));
    defparam mlp_mode_20.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i0 (.D(n62956), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [0]));
    defparam hidden_outputs_0__i0_i0.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i22 (.D(n66298), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [22]));
    defparam output_outputs_1__i0_i22.GSR = "DISABLED";
    FD1P3IX o_4661__i29 (.D(n134_adj_404[29]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[29]));
    defparam o_4661__i29.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i21 (.D(n66454), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [21]));
    defparam output_outputs_1__i0_i21.GSR = "DISABLED";
    FD1P3AX e_i0_i29 (.D(float_alu_c[29]), .SP(n4599), .CK(clock), .Q(e[29]));
    defparam e_i0_i29.GSR = "DISABLED";
    CCU2D n_4659_add_4_13 (.A0(n[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62652), 
          .COUT(n62653), .S0(n134_adj_403[11]), .S1(n134_adj_403[12]));
    defparam n_4659_add_4_13.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_13.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_13.INJECT1_0 = "NO";
    defparam n_4659_add_4_13.INJECT1_1 = "NO";
    FD1P3AX e_i0_i28 (.D(float_alu_c[28]), .SP(n4599), .CK(clock), .Q(e[28]));
    defparam e_i0_i28.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i13 (.D(\hidden_outputs[0] [13]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [13]));
    defparam temp_outputs_0__i0_i13.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i0 (.D(n63188), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [0]));
    defparam hidden_outputs_1__i0_i0.GSR = "DISABLED";
    CCU2D n_4659_add_4_11 (.A0(n[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62651), 
          .COUT(n62652), .S0(n134_adj_403[9]), .S1(n134_adj_403[10]));
    defparam n_4659_add_4_11.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_11.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_11.INJECT1_0 = "NO";
    defparam n_4659_add_4_11.INJECT1_1 = "NO";
    FD1P3IX o_4661__i28 (.D(n134_adj_404[28]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[28]));
    defparam o_4661__i28.GSR = "DISABLED";
    LUT4 i19_4_lut (.A(numL[29]), .B(n38), .C(n28), .D(numL[13]), .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    FD1P3AX output_outputs_1__i0_i20 (.D(n66322), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [20]));
    defparam output_outputs_1__i0_i20.GSR = "DISABLED";
    CCU2D n_4659_add_4_9 (.A0(n[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62650), 
          .COUT(n62651), .S0(n134_adj_403[7]), .S1(n134_adj_403[8]));
    defparam n_4659_add_4_9.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_9.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_9.INJECT1_0 = "NO";
    defparam n_4659_add_4_9.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_7 (.A0(n[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62649), 
          .COUT(n62650), .S0(n134_adj_403[5]), .S1(n134_adj_403[6]));
    defparam n_4659_add_4_7.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_7.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_7.INJECT1_0 = "NO";
    defparam n_4659_add_4_7.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_5 (.A0(n[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62648), 
          .COUT(n62649), .S0(n134_adj_403[3]), .S1(n134_adj_403[4]));
    defparam n_4659_add_4_5.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_5.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_5.INJECT1_0 = "NO";
    defparam n_4659_add_4_5.INJECT1_1 = "NO";
    CCU2D n_4659_add_4_3 (.A0(n[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62647), 
          .COUT(n62648), .S0(n134_adj_403[1]), .S1(n134_adj_403[2]));
    defparam n_4659_add_4_3.INIT0 = 16'hfaaa;
    defparam n_4659_add_4_3.INIT1 = 16'hfaaa;
    defparam n_4659_add_4_3.INJECT1_0 = "NO";
    defparam n_4659_add_4_3.INJECT1_1 = "NO";
    FD1P3IX o_4661__i27 (.D(n134_adj_404[27]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[27]));
    defparam o_4661__i27.GSR = "DISABLED";
    CCU2D n_4659_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62647), 
          .S1(n134_adj_403[0]));
    defparam n_4659_add_4_1.INIT0 = 16'hF000;
    defparam n_4659_add_4_1.INIT1 = 16'h0555;
    defparam n_4659_add_4_1.INJECT1_0 = "NO";
    defparam n_4659_add_4_1.INJECT1_1 = "NO";
    FD1P3AX output_outputs_1__i0_i19 (.D(n66336), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [19]));
    defparam output_outputs_1__i0_i19.GSR = "DISABLED";
    CCU2D o_4661_add_4_33 (.A0(o[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62646), 
          .S0(n134_adj_404[31]));
    defparam o_4661_add_4_33.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_33.INIT1 = 16'h0000;
    defparam o_4661_add_4_33.INJECT1_0 = "NO";
    defparam o_4661_add_4_33.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_31 (.A0(o[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62645), 
          .COUT(n62646), .S0(n134_adj_404[29]), .S1(n134_adj_404[30]));
    defparam o_4661_add_4_31.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_31.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_31.INJECT1_0 = "NO";
    defparam o_4661_add_4_31.INJECT1_1 = "NO";
    FD1P3AX output_outputs_1__i0_i18 (.D(n66338), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [18]));
    defparam output_outputs_1__i0_i18.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i17 (.D(n66456), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [17]));
    defparam output_outputs_1__i0_i17.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i16 (.D(n66334), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [16]));
    defparam output_outputs_1__i0_i16.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i15 (.D(n63246), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [15]));
    defparam output_outputs_1__i0_i15.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i14 (.D(n66458), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [14]));
    defparam output_outputs_1__i0_i14.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i13 (.D(n66460), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [13]));
    defparam output_outputs_1__i0_i13.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i12 (.D(n66390), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [12]));
    defparam output_outputs_1__i0_i12.GSR = "DISABLED";
    CCU2D o_4661_add_4_29 (.A0(o[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62644), 
          .COUT(n62645), .S0(n134_adj_404[27]), .S1(n134_adj_404[28]));
    defparam o_4661_add_4_29.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_29.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_29.INJECT1_0 = "NO";
    defparam o_4661_add_4_29.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_27 (.A0(o[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62643), 
          .COUT(n62644), .S0(n134_adj_404[25]), .S1(n134_adj_404[26]));
    defparam o_4661_add_4_27.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_27.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_27.INJECT1_0 = "NO";
    defparam o_4661_add_4_27.INJECT1_1 = "NO";
    FD1P3AX output_outputs_1__i0_i11 (.D(n66400), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [11]));
    defparam output_outputs_1__i0_i11.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i0 (.D(n66300), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [0]));
    defparam hidden_outputs_2__i0_i0.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i10 (.D(n66526), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [10]));
    defparam output_outputs_1__i0_i10.GSR = "DISABLED";
    FD1P3IX o_4661__i26 (.D(n134_adj_404[26]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[26]));
    defparam o_4661__i26.GSR = "DISABLED";
    CCU2D o_4661_add_4_25 (.A0(o[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62642), 
          .COUT(n62643), .S0(n134_adj_404[23]), .S1(n134_adj_404[24]));
    defparam o_4661_add_4_25.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_25.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_25.INJECT1_0 = "NO";
    defparam o_4661_add_4_25.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_23 (.A0(o[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62641), 
          .COUT(n62642), .S0(n134_adj_404[21]), .S1(n134_adj_404[22]));
    defparam o_4661_add_4_23.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_23.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_23.INJECT1_0 = "NO";
    defparam o_4661_add_4_23.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_0__i0_i2 (.D(\hidden_outputs[0] [2]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [2]));
    defparam temp_outputs_0__i0_i2.GSR = "DISABLED";
    CCU2D o_4661_add_4_21 (.A0(o[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62640), 
          .COUT(n62641), .S0(n134_adj_404[19]), .S1(n134_adj_404[20]));
    defparam o_4661_add_4_21.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_21.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_21.INJECT1_0 = "NO";
    defparam o_4661_add_4_21.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_19 (.A0(o[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62639), 
          .COUT(n62640), .S0(n134_adj_404[17]), .S1(n134_adj_404[18]));
    defparam o_4661_add_4_19.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_19.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_19.INJECT1_0 = "NO";
    defparam o_4661_add_4_19.INJECT1_1 = "NO";
    FD1P3AX e_i0_i27 (.D(float_alu_c[27]), .SP(n4599), .CK(clock), .Q(e[27]));
    defparam e_i0_i27.GSR = "DISABLED";
    FD1P3AX e_i0_i26 (.D(float_alu_c[26]), .SP(n4599), .CK(clock), .Q(e[26]));
    defparam e_i0_i26.GSR = "DISABLED";
    FD1P3AX e_i0_i25 (.D(float_alu_c[25]), .SP(n4599), .CK(clock), .Q(e[25]));
    defparam e_i0_i25.GSR = "DISABLED";
    FD1P3AX e_i0_i24 (.D(float_alu_c[24]), .SP(n4599), .CK(clock), .Q(e[24]));
    defparam e_i0_i24.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n2022[3]), .B(n65), .C(weight_done), .D(n2086), 
         .Z(n2239)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf888;
    CCU2D o_4661_add_4_17 (.A0(o[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62638), 
          .COUT(n62639), .S0(n134_adj_404[15]), .S1(n134_adj_404[16]));
    defparam o_4661_add_4_17.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_17.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_17.INJECT1_0 = "NO";
    defparam o_4661_add_4_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_799_4_lut (.A(n2022[3]), .B(n65), .C(n70822), .D(n2086), 
         .Z(n70769)) /* synthesis lut_function=(A (B (C))+!A (C (D))) */ ;
    defparam i1_4_lut_rep_799_4_lut.init = 16'hd080;
    FD1P3IX o_4661__i25 (.D(n134_adj_404[25]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[25]));
    defparam o_4661__i25.GSR = "DISABLED";
    LUT4 i12333_2_lut_4_lut_3_lut (.A(n2022[3]), .B(n70822), .C(n2086), 
         .Z(n24023)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i12333_2_lut_4_lut_3_lut.init = 16'h4040;
    CCU2D o_4661_add_4_15 (.A0(o[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62637), 
          .COUT(n62638), .S0(n134_adj_404[13]), .S1(n134_adj_404[14]));
    defparam o_4661_add_4_15.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_15.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_15.INJECT1_0 = "NO";
    defparam o_4661_add_4_15.INJECT1_1 = "NO";
    LUT4 i12331_2_lut_3_lut (.A(n2022[27]), .B(n70822), .C(n2086), .Z(n24021)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i12331_2_lut_3_lut.init = 16'h4040;
    CCU2D o_4661_add_4_13 (.A0(o[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62636), 
          .COUT(n62637), .S0(n134_adj_404[11]), .S1(n134_adj_404[12]));
    defparam o_4661_add_4_13.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_13.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_13.INJECT1_0 = "NO";
    defparam o_4661_add_4_13.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_847 (.A(n2022[27]), .B(n70822), .C(n2086), .Z(n70817)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_rep_847.init = 16'hc8c8;
    FD1P3AX output_outputs_1__i0_i9 (.D(n66348), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [9]));
    defparam output_outputs_1__i0_i9.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_2 (.A(n70866), .B(float_alu_ready), .C(n2086), 
         .D(weight_done), .Z(n64)) /* synthesis lut_function=(!(A+!(B ((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_2.init = 16'h4404;
    FD1P3AX output_outputs_1__i0_i8 (.D(n66474), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [8]));
    defparam output_outputs_1__i0_i8.GSR = "DISABLED";
    FD1P3IX o_4661__i24 (.D(n134_adj_404[24]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[24]));
    defparam o_4661__i24.GSR = "DISABLED";
    CCU2D o_4661_add_4_11 (.A0(o[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62635), 
          .COUT(n62636), .S0(n134_adj_404[9]), .S1(n134_adj_404[10]));
    defparam o_4661_add_4_11.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_11.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_11.INJECT1_0 = "NO";
    defparam o_4661_add_4_11.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_9 (.A0(o[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62634), 
          .COUT(n62635), .S0(n134_adj_404[7]), .S1(n134_adj_404[8]));
    defparam o_4661_add_4_9.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_9.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_9.INJECT1_0 = "NO";
    defparam o_4661_add_4_9.INJECT1_1 = "NO";
    FD1P3AX output_outputs_1__i0_i7 (.D(n63058), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [7]));
    defparam output_outputs_1__i0_i7.GSR = "DISABLED";
    CCU2D o_4661_add_4_7 (.A0(o[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62633), 
          .COUT(n62634), .S0(n134_adj_404[5]), .S1(n134_adj_404[6]));
    defparam o_4661_add_4_7.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_7.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_7.INJECT1_0 = "NO";
    defparam o_4661_add_4_7.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_5 (.A0(o[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62632), 
          .COUT(n62633), .S0(n134_adj_404[3]), .S1(n134_adj_404[4]));
    defparam o_4661_add_4_5.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_5.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_5.INJECT1_0 = "NO";
    defparam o_4661_add_4_5.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_3 (.A0(o[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62631), 
          .COUT(n62632), .S0(n134_adj_404[1]), .S1(n134_adj_404[2]));
    defparam o_4661_add_4_3.INIT0 = 16'hfaaa;
    defparam o_4661_add_4_3.INIT1 = 16'hfaaa;
    defparam o_4661_add_4_3.INJECT1_0 = "NO";
    defparam o_4661_add_4_3.INJECT1_1 = "NO";
    CCU2D o_4661_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62631), 
          .S1(n134_adj_404[0]));
    defparam o_4661_add_4_1.INIT0 = 16'hF000;
    defparam o_4661_add_4_1.INIT1 = 16'h0555;
    defparam o_4661_add_4_1.INJECT1_0 = "NO";
    defparam o_4661_add_4_1.INJECT1_1 = "NO";
    FD1P3AX hidden_outputs_3__i0_i0 (.D(n66386), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [0]));
    defparam hidden_outputs_3__i0_i0.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i1 (.D(\hidden_outputs[0] [1]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [1]));
    defparam temp_outputs_0__i0_i1.GSR = "DISABLED";
    FD1P3AX e_i0_i23 (.D(float_alu_c[23]), .SP(n4599), .CK(clock), .Q(e[23]));
    defparam e_i0_i23.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i0 (.D(n63022), .SP(n23664), .CK(clock), .Q(float_alu_b[0]));
    defparam float_alu_b_i0_i0.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i6 (.D(n66292), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [6]));
    defparam output_outputs_1__i0_i6.GSR = "DISABLED";
    FD1P3IX o_4661__i23 (.D(n134_adj_404[23]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[23]));
    defparam o_4661__i23.GSR = "DISABLED";
    DPR16X4C inputs6 (.DI0(sram_output_B[4]), .DI1(sram_output_B[5]), .DI2(sram_output_B[6]), 
            .DI3(sram_output_B[7]), .WAD0(addr[0]), .WAD1(addr[1]), .WAD2(addr[2]), 
            .WAD3(GND_net), .WCK(clock), .WRE(n15113), .RAD0(i[0]), 
            .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), .DO0(n1027[4]), 
            .DO1(n1027[5]), .DO2(n1027[6]), .DO3(n1027[7]));
    defparam inputs6.initval = "0x0000000000000000";
    FD1P3AX temp_outputs_1__i0_i31 (.D(\hidden_outputs[1] [31]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [31]));
    defparam temp_outputs_1__i0_i31.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i30 (.D(\hidden_outputs[1] [30]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [30]));
    defparam temp_outputs_1__i0_i30.GSR = "DISABLED";
    DPR16X4C inputs5 (.DI0(sram_output_B[8]), .DI1(sram_output_B[9]), .DI2(sram_output_B[10]), 
            .DI3(sram_output_B[11]), .WAD0(addr[0]), .WAD1(addr[1]), .WAD2(addr[2]), 
            .WAD3(GND_net), .WCK(clock), .WRE(n15113), .RAD0(i[0]), 
            .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), .DO0(n1027[8]), 
            .DO1(n1027[9]), .DO2(n1027[10]), .DO3(n1027[11]));
    defparam inputs5.initval = "0x0000000000000000";
    DPR16X4C inputs4 (.DI0(sram_output_B[12]), .DI1(sram_output_B[13]), 
            .DI2(sram_output_B[14]), .DI3(sram_output_B[15]), .WAD0(addr[0]), 
            .WAD1(addr[1]), .WAD2(addr[2]), .WAD3(GND_net), .WCK(clock), 
            .WRE(n15113), .RAD0(i[0]), .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), 
            .DO0(n1027[12]), .DO1(n1027[13]), .DO2(n1027[14]), .DO3(n1027[15]));
    defparam inputs4.initval = "0x0000000000000000";
    FD1P3AX output_outputs_1__i0_i5 (.D(n66468), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [5]));
    defparam output_outputs_1__i0_i5.GSR = "DISABLED";
    DPR16X4C inputs3 (.DI0(sram_output_B[16]), .DI1(sram_output_B[17]), 
            .DI2(sram_output_B[18]), .DI3(sram_output_B[19]), .WAD0(addr[0]), 
            .WAD1(addr[1]), .WAD2(addr[2]), .WAD3(GND_net), .WCK(clock), 
            .WRE(n15113), .RAD0(i[0]), .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), 
            .DO0(n1027[16]), .DO1(n1027[17]), .DO2(n1027[18]), .DO3(n1027[19]));
    defparam inputs3.initval = "0x0000000000000000";
    FD1P3AX e_i0_i22 (.D(float_alu_c[22]), .SP(n4599), .CK(clock), .Q(e[22]));
    defparam e_i0_i22.GSR = "DISABLED";
    FD1P3AX e_i0_i21 (.D(float_alu_c[21]), .SP(n4599), .CK(clock), .Q(e[21]));
    defparam e_i0_i21.GSR = "DISABLED";
    FD1P3AX e_i0_i20 (.D(float_alu_c[20]), .SP(n4599), .CK(clock), .Q(e[20]));
    defparam e_i0_i20.GSR = "DISABLED";
    FD1P3AX e_i0_i19 (.D(float_alu_c[19]), .SP(n4599), .CK(clock), .Q(e[19]));
    defparam e_i0_i19.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i0 (.D(n66466), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [0]));
    defparam hidden_outputs_4__i0_i0.GSR = "DISABLED";
    CCU2D add_4584_add_1_add_1_7 (.A0(n14054), .B0(numL[0]), .C0(n12), 
          .D0(n927), .A1(n14054), .B1(numL[0]), .C1(n12), .D1(n926), 
          .CIN(n61484), .COUT(n61485), .S0(n3[5]), .S1(n3[6]));
    defparam add_4584_add_1_add_1_7.INIT0 = 16'hfe00;
    defparam add_4584_add_1_add_1_7.INIT1 = 16'hfe00;
    defparam add_4584_add_1_add_1_7.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_7.INJECT1_1 = "NO";
    FD1P3AX e_i0_i18 (.D(float_alu_c[18]), .SP(n4599), .CK(clock), .Q(e[18]));
    defparam e_i0_i18.GSR = "DISABLED";
    FD1P3AX e_i0_i17 (.D(float_alu_c[17]), .SP(n4599), .CK(clock), .Q(e[17]));
    defparam e_i0_i17.GSR = "DISABLED";
    FD1P3AX e_i0_i16 (.D(float_alu_c[16]), .SP(n4599), .CK(clock), .Q(e[16]));
    defparam e_i0_i16.GSR = "DISABLED";
    FD1P3AX e_i0_i15 (.D(float_alu_c[15]), .SP(n4599), .CK(clock), .Q(e[15]));
    defparam e_i0_i15.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i4 (.D(n63047), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [4]));
    defparam output_outputs_1__i0_i4.GSR = "DISABLED";
    FD1P3AX e_i0_i14 (.D(float_alu_c[14]), .SP(n4599), .CK(clock), .Q(e[14]));
    defparam e_i0_i14.GSR = "DISABLED";
    DPR16X4C inputs2 (.DI0(sram_output_B[20]), .DI1(sram_output_B[21]), 
            .DI2(sram_output_B[22]), .DI3(sram_output_B[23]), .WAD0(addr[0]), 
            .WAD1(addr[1]), .WAD2(addr[2]), .WAD3(GND_net), .WCK(clock), 
            .WRE(n15113), .RAD0(i[0]), .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), 
            .DO0(n1027[20]), .DO1(n1027[21]), .DO2(n1027[22]), .DO3(n1027[23]));
    defparam inputs2.initval = "0x0000000000000000";
    FD1P3AX e_i0_i13 (.D(float_alu_c[13]), .SP(n4599), .CK(clock), .Q(e[13]));
    defparam e_i0_i13.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i3 (.D(n66530), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [3]));
    defparam output_outputs_1__i0_i3.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i2 (.D(n66306), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [2]));
    defparam output_outputs_1__i0_i2.GSR = "DISABLED";
    FD1P3AX output_outputs_1__i0_i1 (.D(n63077), .SP(n23647), .CK(clock), 
            .Q(\mlp_outputs[1] [1]));
    defparam output_outputs_1__i0_i1.GSR = "DISABLED";
    FD1P3IX o_4661__i22 (.D(n134_adj_404[22]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[22]));
    defparam o_4661__i22.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(float_alu_ready), .B(n70866), .C(SDA_c), .D(n2022[28]), 
         .Z(n4613)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0200;
    FD1P3IX o_4661__i21 (.D(n134_adj_404[21]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[21]));
    defparam o_4661__i21.GSR = "DISABLED";
    FD1P3AX temp_outputs_1__i0_i29 (.D(\hidden_outputs[1] [29]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [29]));
    defparam temp_outputs_1__i0_i29.GSR = "DISABLED";
    FD1P3AX e_i0_i12 (.D(float_alu_c[12]), .SP(n4599), .CK(clock), .Q(e[12]));
    defparam e_i0_i12.GSR = "DISABLED";
    CCU2D counter_4663_4767_add_4_13 (.A0(counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62613), .S0(n54[11]));
    defparam counter_4663_4767_add_4_13.INIT0 = 16'hfaaa;
    defparam counter_4663_4767_add_4_13.INIT1 = 16'h0000;
    defparam counter_4663_4767_add_4_13.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_13.INJECT1_1 = "NO";
    FD1P3AX e_i0_i11 (.D(float_alu_c[11]), .SP(n4599), .CK(clock), .Q(e[11]));
    defparam e_i0_i11.GSR = "DISABLED";
    CCU2D counter_4663_4767_add_4_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62612), .COUT(n62613), .S0(n54[9]), .S1(n54[10]));
    defparam counter_4663_4767_add_4_11.INIT0 = 16'hfaaa;
    defparam counter_4663_4767_add_4_11.INIT1 = 16'hfaaa;
    defparam counter_4663_4767_add_4_11.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_11.INJECT1_1 = "NO";
    FD1P3DX ready_78 (.D(n70788), .SP(n70778), .CK(clock), .CD(SDA_c), 
            .Q(float_alu_ready));
    defparam ready_78.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_rep_909 (.A(n70731), .B(n14054), .C(n4613), 
         .D(numL[31]), .Z(n73807)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_rep_909.init = 16'hf010;
    DPR16X4C inputs7 (.DI0(sram_output_B[0]), .DI1(sram_output_B[1]), .DI2(sram_output_B[2]), 
            .DI3(sram_output_B[3]), .WAD0(addr[0]), .WAD1(addr[1]), .WAD2(addr[2]), 
            .WAD3(GND_net), .WCK(clock), .WRE(n15113), .RAD0(i[0]), 
            .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), .DO0(n1027[0]), 
            .DO1(n1027[1]), .DO2(n1027[2]), .DO3(n1027[3]));
    defparam inputs7.initval = "0x0000000000000000";
    LUT4 i6567_1_lut (.A(n14054), .Z(n14050)) /* synthesis lut_function=(!(A)) */ ;
    defparam i6567_1_lut.init = 16'h5555;
    FD1P3IX o_4661__i20 (.D(n134_adj_404[20]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[20]));
    defparam o_4661__i20.GSR = "DISABLED";
    CCU2D counter_4663_4767_add_4_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62611), .COUT(n62612), .S0(n54[7]), .S1(n54[8]));
    defparam counter_4663_4767_add_4_9.INIT0 = 16'hfaaa;
    defparam counter_4663_4767_add_4_9.INIT1 = 16'hfaaa;
    defparam counter_4663_4767_add_4_9.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_9.INJECT1_1 = "NO";
    FD1P3IX o_4661__i19 (.D(n134_adj_404[19]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[19]));
    defparam o_4661__i19.GSR = "DISABLED";
    CCU2D counter_4663_4767_add_4_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n62610), .COUT(n62611), .S0(n54[5]), .S1(n54[6]));
    defparam counter_4663_4767_add_4_7.INIT0 = 16'hfaaa;
    defparam counter_4663_4767_add_4_7.INIT1 = 16'hfaaa;
    defparam counter_4663_4767_add_4_7.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_7.INJECT1_1 = "NO";
    CCU2D equal_97_28 (.A0(i_c[19]), .B0(i_c[18]), .C0(i_c[17]), .D0(i_c[16]), 
          .A1(i_c[16]), .B1(i_c[15]), .C1(i_c[14]), .D1(i_c[13]), .CIN(n60975), 
          .COUT(n60976));
    defparam equal_97_28.INIT0 = 16'h8001;
    defparam equal_97_28.INIT1 = 16'h8001;
    defparam equal_97_28.INJECT1_0 = "YES";
    defparam equal_97_28.INJECT1_1 = "YES";
    FD1P3AX e_i0_i10 (.D(float_alu_c[10]), .SP(n4599), .CK(clock), .Q(e[10]));
    defparam e_i0_i10.GSR = "DISABLED";
    CCU2D equal_97_26 (.A0(i_c[25]), .B0(i_c[24]), .C0(i_c[23]), .D0(i_c[22]), 
          .A1(i_c[22]), .B1(i_c[21]), .C1(i_c[20]), .D1(i_c[19]), .CIN(n60974), 
          .COUT(n60975));
    defparam equal_97_26.INIT0 = 16'h8001;
    defparam equal_97_26.INIT1 = 16'h8001;
    defparam equal_97_26.INJECT1_0 = "YES";
    defparam equal_97_26.INJECT1_1 = "YES";
    FD1P3AX e_i0_i9 (.D(float_alu_c[9]), .SP(n4599), .CK(clock), .Q(e[9]));
    defparam e_i0_i9.GSR = "DISABLED";
    FD1P3AX e_i0_i8 (.D(float_alu_c[8]), .SP(n4599), .CK(clock), .Q(e[8]));
    defparam e_i0_i8.GSR = "DISABLED";
    FD1P3AX e_i0_i7 (.D(float_alu_c[7]), .SP(n4599), .CK(clock), .Q(e[7]));
    defparam e_i0_i7.GSR = "DISABLED";
    CCU2D counter_4663_4767_add_4_5 (.A0(counter[3]), .B0(n70713), .C0(n2889[3]), 
          .D0(n3044[3]), .A1(counter[4]), .B1(n70713), .C1(n2889[4]), 
          .D1(n3044[4]), .CIN(n62609), .COUT(n62610), .S0(n54[3]), .S1(n54[4]));
    defparam counter_4663_4767_add_4_5.INIT0 = 16'h596a;
    defparam counter_4663_4767_add_4_5.INIT1 = 16'h596a;
    defparam counter_4663_4767_add_4_5.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_5.INJECT1_1 = "NO";
    FD1P3IX o_4661__i18 (.D(n134_adj_404[18]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[18]));
    defparam o_4661__i18.GSR = "DISABLED";
    CCU2D counter_4663_4767_add_4_3 (.A0(counter[1]), .B0(n70713), .C0(n2889[1]), 
          .D0(n3044[1]), .A1(counter[2]), .B1(n70713), .C1(n2889[2]), 
          .D1(n3044[2]), .CIN(n62608), .COUT(n62609), .S0(n54[1]), .S1(n54[2]));
    defparam counter_4663_4767_add_4_3.INIT0 = 16'h596a;
    defparam counter_4663_4767_add_4_3.INIT1 = 16'h596a;
    defparam counter_4663_4767_add_4_3.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_3.INJECT1_1 = "NO";
    CCU2D counter_4663_4767_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[0]), .B1(n70713), .C1(n2889[0]), 
          .D1(n3044[0]), .COUT(n62608), .S1(n54[0]));
    defparam counter_4663_4767_add_4_1.INIT0 = 16'hF000;
    defparam counter_4663_4767_add_4_1.INIT1 = 16'h596a;
    defparam counter_4663_4767_add_4_1.INJECT1_0 = "NO";
    defparam counter_4663_4767_add_4_1.INJECT1_1 = "NO";
    FD1P3AX e_i0_i6 (.D(float_alu_c[6]), .SP(n4599), .CK(clock), .Q(e[6]));
    defparam e_i0_i6.GSR = "DISABLED";
    CCU2D add_4994_11 (.A0(h[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62606), 
          .S0(n7702[9]), .S1(n7702[10]));
    defparam add_4994_11.INIT0 = 16'hfaaa;
    defparam add_4994_11.INIT1 = 16'hfaaa;
    defparam add_4994_11.INJECT1_0 = "NO";
    defparam add_4994_11.INJECT1_1 = "NO";
    CCU2D add_4994_9 (.A0(h[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62605), 
          .COUT(n62606), .S0(n7702[7]), .S1(n7702[8]));
    defparam add_4994_9.INIT0 = 16'hfaaa;
    defparam add_4994_9.INIT1 = 16'hfaaa;
    defparam add_4994_9.INJECT1_0 = "NO";
    defparam add_4994_9.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_0__i0_i12 (.D(\hidden_outputs[0] [12]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [12]));
    defparam temp_outputs_0__i0_i12.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i11 (.D(\hidden_outputs[0] [11]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [11]));
    defparam temp_outputs_0__i0_i11.GSR = "DISABLED";
    DPR16X4C inputs0 (.DI0(sram_output_B[28]), .DI1(sram_output_B[29]), 
            .DI2(sram_output_B[30]), .DI3(sram_output_B[31]), .WAD0(addr[0]), 
            .WAD1(addr[1]), .WAD2(addr[2]), .WAD3(GND_net), .WCK(clock), 
            .WRE(n15113), .RAD0(i[0]), .RAD1(i[1]), .RAD2(i[2]), .RAD3(GND_net), 
            .DO0(n1027[28]), .DO1(n1027[29]), .DO2(n1027[30]), .DO3(n1027[31]));
    defparam inputs0.initval = "0x0000000000000000";
    FD1P3AX e_i0_i5 (.D(float_alu_c[5]), .SP(n4599), .CK(clock), .Q(e[5]));
    defparam e_i0_i5.GSR = "DISABLED";
    CCU2D add_4994_7 (.A0(h[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62604), 
          .COUT(n62605), .S0(n7702[5]), .S1(n7702[6]));
    defparam add_4994_7.INIT0 = 16'hfaaa;
    defparam add_4994_7.INIT1 = 16'hfaaa;
    defparam add_4994_7.INJECT1_0 = "NO";
    defparam add_4994_7.INJECT1_1 = "NO";
    CCU2D add_4994_5 (.A0(h[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62603), 
          .COUT(n62604), .S0(n7702[3]), .S1(n7702[4]));
    defparam add_4994_5.INIT0 = 16'hfaaa;
    defparam add_4994_5.INIT1 = 16'hfaaa;
    defparam add_4994_5.INJECT1_0 = "NO";
    defparam add_4994_5.INJECT1_1 = "NO";
    FD1P3AX e_i0_i4 (.D(float_alu_c[4]), .SP(n4599), .CK(clock), .Q(e[4]));
    defparam e_i0_i4.GSR = "DISABLED";
    CCU2D add_4994_3 (.A0(h[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62602), 
          .COUT(n62603), .S0(n7702[1]), .S1(n7702[2]));
    defparam add_4994_3.INIT0 = 16'hfaaa;
    defparam add_4994_3.INIT1 = 16'h0555;
    defparam add_4994_3.INJECT1_0 = "NO";
    defparam add_4994_3.INJECT1_1 = "NO";
    FD1P3AX e_i0_i3 (.D(float_alu_c[3]), .SP(n4599), .CK(clock), .Q(e[3]));
    defparam e_i0_i3.GSR = "DISABLED";
    FD1P3AX e_i0_i2 (.D(float_alu_c[2]), .SP(n4599), .CK(clock), .Q(e[2]));
    defparam e_i0_i2.GSR = "DISABLED";
    LUT4 i9_2_lut (.A(numL[20]), .B(numL[8]), .Z(n32)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    FD1P3AX e_i0_i1 (.D(float_alu_c[1]), .SP(n4599), .CK(clock), .Q(e[1]));
    defparam e_i0_i1.GSR = "DISABLED";
    FD1P3AX weight_i0_i31 (.D(sram_output_B[31]), .SP(n4593), .CK(clock), 
            .Q(weight[31]));
    defparam weight_i0_i31.GSR = "DISABLED";
    FD1P3AX weight_i0_i30 (.D(sram_output_B[30]), .SP(n4593), .CK(clock), 
            .Q(weight[30]));
    defparam weight_i0_i30.GSR = "DISABLED";
    FD1P3AX weight_i0_i29 (.D(sram_output_B[29]), .SP(n4593), .CK(clock), 
            .Q(weight[29]));
    defparam weight_i0_i29.GSR = "DISABLED";
    FD1P3AX weight_i0_i28 (.D(sram_output_B[28]), .SP(n4593), .CK(clock), 
            .Q(weight[28]));
    defparam weight_i0_i28.GSR = "DISABLED";
    FD1P3AX weight_i0_i27 (.D(sram_output_B[27]), .SP(n4593), .CK(clock), 
            .Q(weight[27]));
    defparam weight_i0_i27.GSR = "DISABLED";
    FD1P3AX weight_i0_i26 (.D(sram_output_B[26]), .SP(n4593), .CK(clock), 
            .Q(weight[26]));
    defparam weight_i0_i26.GSR = "DISABLED";
    FD1P3AX weight_i0_i25 (.D(sram_output_B[25]), .SP(n4593), .CK(clock), 
            .Q(weight[25]));
    defparam weight_i0_i25.GSR = "DISABLED";
    FD1P3AX weight_i0_i24 (.D(sram_output_B[24]), .SP(n4593), .CK(clock), 
            .Q(weight[24]));
    defparam weight_i0_i24.GSR = "DISABLED";
    FD1P3AX weight_i0_i23 (.D(sram_output_B[23]), .SP(n4593), .CK(clock), 
            .Q(weight[23]));
    defparam weight_i0_i23.GSR = "DISABLED";
    FD1P3AX weight_i0_i22 (.D(sram_output_B[22]), .SP(n4593), .CK(clock), 
            .Q(weight[22]));
    defparam weight_i0_i22.GSR = "DISABLED";
    FD1P3AX weight_i0_i21 (.D(sram_output_B[21]), .SP(n4593), .CK(clock), 
            .Q(weight[21]));
    defparam weight_i0_i21.GSR = "DISABLED";
    FD1P3AX weight_i0_i20 (.D(sram_output_B[20]), .SP(n4593), .CK(clock), 
            .Q(weight[20]));
    defparam weight_i0_i20.GSR = "DISABLED";
    FD1P3AX weight_i0_i19 (.D(sram_output_B[19]), .SP(n4593), .CK(clock), 
            .Q(weight[19]));
    defparam weight_i0_i19.GSR = "DISABLED";
    FD1P3AX weight_i0_i18 (.D(sram_output_B[18]), .SP(n4593), .CK(clock), 
            .Q(weight[18]));
    defparam weight_i0_i18.GSR = "DISABLED";
    FD1P3AX weight_i0_i17 (.D(sram_output_B[17]), .SP(n4593), .CK(clock), 
            .Q(weight[17]));
    defparam weight_i0_i17.GSR = "DISABLED";
    FD1P3AX weight_i0_i16 (.D(sram_output_B[16]), .SP(n4593), .CK(clock), 
            .Q(weight[16]));
    defparam weight_i0_i16.GSR = "DISABLED";
    FD1P3AX weight_i0_i15 (.D(sram_output_B[15]), .SP(n4593), .CK(clock), 
            .Q(weight[15]));
    defparam weight_i0_i15.GSR = "DISABLED";
    FD1P3AX weight_i0_i14 (.D(sram_output_B[14]), .SP(n4593), .CK(clock), 
            .Q(weight[14]));
    defparam weight_i0_i14.GSR = "DISABLED";
    FD1P3AX weight_i0_i13 (.D(sram_output_B[13]), .SP(n4593), .CK(clock), 
            .Q(weight[13]));
    defparam weight_i0_i13.GSR = "DISABLED";
    FD1P3AX weight_i0_i12 (.D(sram_output_B[12]), .SP(n4593), .CK(clock), 
            .Q(weight[12]));
    defparam weight_i0_i12.GSR = "DISABLED";
    FD1P3AX weight_i0_i11 (.D(sram_output_B[11]), .SP(n4593), .CK(clock), 
            .Q(weight[11]));
    defparam weight_i0_i11.GSR = "DISABLED";
    FD1P3AX weight_i0_i10 (.D(sram_output_B[10]), .SP(n4593), .CK(clock), 
            .Q(weight[10]));
    defparam weight_i0_i10.GSR = "DISABLED";
    FD1P3AX weight_i0_i9 (.D(sram_output_B[9]), .SP(n4593), .CK(clock), 
            .Q(weight[9]));
    defparam weight_i0_i9.GSR = "DISABLED";
    FD1P3AX weight_i0_i8 (.D(sram_output_B[8]), .SP(n4593), .CK(clock), 
            .Q(weight[8]));
    defparam weight_i0_i8.GSR = "DISABLED";
    FD1P3AX weight_i0_i7 (.D(sram_output_B[7]), .SP(n4593), .CK(clock), 
            .Q(weight[7]));
    defparam weight_i0_i7.GSR = "DISABLED";
    FD1P3AX weight_i0_i6 (.D(sram_output_B[6]), .SP(n4593), .CK(clock), 
            .Q(weight[6]));
    defparam weight_i0_i6.GSR = "DISABLED";
    FD1P3AX weight_i0_i5 (.D(sram_output_B[5]), .SP(n4593), .CK(clock), 
            .Q(weight[5]));
    defparam weight_i0_i5.GSR = "DISABLED";
    FD1P3AX weight_i0_i4 (.D(sram_output_B[4]), .SP(n4593), .CK(clock), 
            .Q(weight[4]));
    defparam weight_i0_i4.GSR = "DISABLED";
    FD1P3AX weight_i0_i3 (.D(sram_output_B[3]), .SP(n4593), .CK(clock), 
            .Q(weight[3]));
    defparam weight_i0_i3.GSR = "DISABLED";
    FD1P3AX weight_i0_i2 (.D(sram_output_B[2]), .SP(n4593), .CK(clock), 
            .Q(weight[2]));
    defparam weight_i0_i2.GSR = "DISABLED";
    FD1P3AX weight_i0_i1 (.D(sram_output_B[1]), .SP(n4593), .CK(clock), 
            .Q(weight[1]));
    defparam weight_i0_i1.GSR = "DISABLED";
    FD1P3IX o_4661__i17 (.D(n134_adj_404[17]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[17]));
    defparam o_4661__i17.GSR = "DISABLED";
    CCU2D add_4994_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62602), 
          .S1(n7702[0]));
    defparam add_4994_1.INIT0 = 16'hF000;
    defparam add_4994_1.INIT1 = 16'h0555;
    defparam add_4994_1.INJECT1_0 = "NO";
    defparam add_4994_1.INJECT1_1 = "NO";
    CCU2D add_49686_12 (.A0(n3_adj_405[10]), .B0(n3_adj_406[10]), .C0(GND_net), 
          .D0(GND_net), .A1(n3_adj_405[11]), .B1(n3_adj_406[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62600), .S0(n61312[10]), .S1(n61312[11]));
    defparam add_49686_12.INIT0 = 16'h5666;
    defparam add_49686_12.INIT1 = 16'h5666;
    defparam add_49686_12.INJECT1_0 = "NO";
    defparam add_49686_12.INJECT1_1 = "NO";
    FD1P3IX o_4661__i16 (.D(n134_adj_404[16]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[16]));
    defparam o_4661__i16.GSR = "DISABLED";
    FD1P3IX o_4661__i15 (.D(n134_adj_404[15]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[15]));
    defparam o_4661__i15.GSR = "DISABLED";
    CCU2D add_49686_10 (.A0(n3_adj_405[8]), .B0(n3_adj_406[8]), .C0(GND_net), 
          .D0(GND_net), .A1(n3_adj_405[9]), .B1(n3_adj_406[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62599), .COUT(n62600), .S0(n61312[8]), 
          .S1(n61312[9]));
    defparam add_49686_10.INIT0 = 16'h5666;
    defparam add_49686_10.INIT1 = 16'h5666;
    defparam add_49686_10.INJECT1_0 = "NO";
    defparam add_49686_10.INJECT1_1 = "NO";
    CCU2D add_49686_8 (.A0(n3_adj_405[6]), .B0(n3_adj_406[6]), .C0(GND_net), 
          .D0(GND_net), .A1(n3_adj_405[7]), .B1(n3_adj_406[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62598), .COUT(n62599), .S0(n61312[6]), 
          .S1(n61312[7]));
    defparam add_49686_8.INIT0 = 16'h5666;
    defparam add_49686_8.INIT1 = 16'h5666;
    defparam add_49686_8.INJECT1_0 = "NO";
    defparam add_49686_8.INJECT1_1 = "NO";
    LUT4 i17_4_lut (.A(numL[27]), .B(numL[14]), .C(numL[4]), .D(numL[21]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    CCU2D add_49686_6 (.A0(n3_adj_405[4]), .B0(n3_adj_406[4]), .C0(GND_net), 
          .D0(GND_net), .A1(n3_adj_405[5]), .B1(n3_adj_406[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62597), .COUT(n62598), .S0(n61312[4]), 
          .S1(n61312[5]));
    defparam add_49686_6.INIT0 = 16'h5666;
    defparam add_49686_6.INIT1 = 16'h5666;
    defparam add_49686_6.INJECT1_0 = "NO";
    defparam add_49686_6.INJECT1_1 = "NO";
    CCU2D add_49686_4 (.A0(n3_adj_405[2]), .B0(n3_adj_406[2]), .C0(GND_net), 
          .D0(GND_net), .A1(n3_adj_405[3]), .B1(n3_adj_406[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n62596), .COUT(n62597), .S0(n61312[2]), 
          .S1(n61312[3]));
    defparam add_49686_4.INIT0 = 16'h5666;
    defparam add_49686_4.INIT1 = 16'h5666;
    defparam add_49686_4.INJECT1_0 = "NO";
    defparam add_49686_4.INJECT1_1 = "NO";
    CCU2D add_49686_2 (.A0(n3_adj_405[0]), .B0(counter[0]), .C0(GND_net), 
          .D0(GND_net), .A1(counter[1]), .B1(n[0]), .C1(n3_adj_405[1]), 
          .D1(GND_net), .COUT(n62596), .S1(n61312[1]));
    defparam add_49686_2.INIT0 = 16'h7000;
    defparam add_49686_2.INIT1 = 16'h9696;
    defparam add_49686_2.INJECT1_0 = "NO";
    defparam add_49686_2.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_798_4_lut (.A(n70860), .B(n70863), .C(n128), .D(n70857), 
         .Z(n70768)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_798_4_lut.init = 16'hfffe;
    CCU2D add_49684_13 (.A0(n12), .B0(n5), .C0(h[11]), .D0(n7702[10]), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62594), 
          .S0(n61292[11]));
    defparam add_49684_13.INIT0 = 16'hf1e0;
    defparam add_49684_13.INIT1 = 16'h0000;
    defparam add_49684_13.INJECT1_0 = "NO";
    defparam add_49684_13.INJECT1_1 = "NO";
    CCU2D add_49684_11 (.A0(n12), .B0(n5), .C0(h[9]), .D0(n7702[8]), 
          .A1(n12), .B1(n5), .C1(h[10]), .D1(n7702[9]), .CIN(n62593), 
          .COUT(n62594), .S0(n61292[9]), .S1(n61292[10]));
    defparam add_49684_11.INIT0 = 16'hf1e0;
    defparam add_49684_11.INIT1 = 16'hf1e0;
    defparam add_49684_11.INJECT1_0 = "NO";
    defparam add_49684_11.INJECT1_1 = "NO";
    FD1P3IX o_4661__i14 (.D(n134_adj_404[14]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[14]));
    defparam o_4661__i14.GSR = "DISABLED";
    CCU2D add_49684_9 (.A0(n12), .B0(n5), .C0(h[7]), .D0(n7702[6]), 
          .A1(n12), .B1(n5), .C1(h[8]), .D1(n7702[7]), .CIN(n62592), 
          .COUT(n62593), .S0(n61292[7]), .S1(n61292[8]));
    defparam add_49684_9.INIT0 = 16'hf1e0;
    defparam add_49684_9.INIT1 = 16'hf1e0;
    defparam add_49684_9.INJECT1_0 = "NO";
    defparam add_49684_9.INJECT1_1 = "NO";
    CCU2D add_49684_7 (.A0(n12), .B0(n5), .C0(h[5]), .D0(n7702[4]), 
          .A1(n12), .B1(n5), .C1(h[6]), .D1(n7702[5]), .CIN(n62591), 
          .COUT(n62592), .S0(n61292[5]), .S1(n61292[6]));
    defparam add_49684_7.INIT0 = 16'hf1e0;
    defparam add_49684_7.INIT1 = 16'hf1e0;
    defparam add_49684_7.INJECT1_0 = "NO";
    defparam add_49684_7.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i28 (.D(\hidden_outputs[1] [28]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [28]));
    defparam temp_outputs_1__i0_i28.GSR = "DISABLED";
    CCU2D add_49684_5 (.A0(n66817), .B0(n70712), .C0(h[3]), .D0(n7702[2]), 
          .A1(n13918[4]), .B1(n66247), .C1(n65435), .D1(n15041[3]), 
          .CIN(n62590), .COUT(n62591), .S0(n61292[3]), .S1(n61292[4]));
    defparam add_49684_5.INIT0 = 16'h596a;
    defparam add_49684_5.INIT1 = 16'h56aa;
    defparam add_49684_5.INJECT1_0 = "NO";
    defparam add_49684_5.INJECT1_1 = "NO";
    CCU2D add_49684_3 (.A0(n70712), .B0(n61391), .C0(h[1]), .D0(n7702[0]), 
          .A1(n13918[2]), .B1(n70712), .C1(n70708), .D1(n236[2]), .CIN(n62589), 
          .COUT(n62590), .S0(n61292[1]), .S1(n61292[2]));
    defparam add_49684_3.INIT0 = 16'h7d28;
    defparam add_49684_3.INIT1 = 16'h5a96;
    defparam add_49684_3.INJECT1_0 = "NO";
    defparam add_49684_3.INJECT1_1 = "NO";
    CCU2D add_49684_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(h[0]), .B1(n12), .C1(n5), .D1(n61382), .COUT(n62589), 
          .S1(n61292[0]));
    defparam add_49684_1.INIT0 = 16'hF000;
    defparam add_49684_1.INIT1 = 16'h56aa;
    defparam add_49684_1.INJECT1_0 = "NO";
    defparam add_49684_1.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i27 (.D(\hidden_outputs[1] [27]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [27]));
    defparam temp_outputs_1__i0_i27.GSR = "DISABLED";
    CCU2D add_49683_13 (.A0(n61292[11]), .B0(n12), .C0(n5), .D0(counter[11]), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62588), 
          .S0(n61278[11]));
    defparam add_49683_13.INIT0 = 16'h56aa;
    defparam add_49683_13.INIT1 = 16'h0000;
    defparam add_49683_13.INJECT1_0 = "NO";
    defparam add_49683_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_3 (.A(n2022[38]), .B(n10_adj_71), .C(n2022[45]), 
         .D(n2022[39]), .Z(n4_adj_72)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_3.init = 16'hfffe;
    LUT4 i5_3_lut_rep_839 (.A(n2022[38]), .B(n10_adj_71), .C(n2022[45]), 
         .Z(n70809)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut_rep_839.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_4 (.A(n2022[31]), .B(n70822), .C(n46466), 
         .D(o[0]), .Z(n23647)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut_adj_4.init = 16'hf8f0;
    LUT4 i1_3_lut_4_lut_adj_5 (.A(n2022[31]), .B(n70822), .C(n46466), 
         .D(o[0]), .Z(n23646)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;
    defparam i1_3_lut_4_lut_adj_5.init = 16'hf0f8;
    CCU2D add_49683_11 (.A0(n61292[9]), .B0(n12), .C0(n5), .D0(counter[9]), 
          .A1(n61292[10]), .B1(n12), .C1(n5), .D1(counter[10]), .CIN(n62587), 
          .COUT(n62588), .S0(n61278[9]), .S1(n61278[10]));
    defparam add_49683_11.INIT0 = 16'h56aa;
    defparam add_49683_11.INIT1 = 16'h56aa;
    defparam add_49683_11.INJECT1_0 = "NO";
    defparam add_49683_11.INJECT1_1 = "NO";
    LUT4 select_455_Select_1_i32_2_lut (.A(sram_output_B[1]), .B(n2022[31]), 
         .Z(n32_adj_73)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_1_i32_2_lut.init = 16'h8888;
    CCU2D add_49683_9 (.A0(n61292[7]), .B0(n12), .C0(n5), .D0(counter[7]), 
          .A1(n61292[8]), .B1(n12), .C1(n5), .D1(counter[8]), .CIN(n62586), 
          .COUT(n62587), .S0(n61278[7]), .S1(n61278[8]));
    defparam add_49683_9.INIT0 = 16'h56aa;
    defparam add_49683_9.INIT1 = 16'h56aa;
    defparam add_49683_9.INJECT1_0 = "NO";
    defparam add_49683_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(\mlp_outputs[1] [1]), .B(n70809), .C(float_alu_c[1]), 
         .D(o[0]), .Z(n23234)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i2_4_lut (.A(n23234), .B(n32_adj_73), .C(\mlp_outputs[1] [1]), 
         .D(n2022[39]), .Z(n63077)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'hfeee;
    LUT4 i21_4_lut (.A(numL[9]), .B(n42), .C(n36), .D(n24), .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    CCU2D add_49683_7 (.A0(n61292[5]), .B0(n12), .C0(n5), .D0(counter[5]), 
          .A1(n61292[6]), .B1(n12), .C1(n5), .D1(counter[6]), .CIN(n62585), 
          .COUT(n62586), .S0(n61278[5]), .S1(n61278[6]));
    defparam add_49683_7.INIT0 = 16'h56aa;
    defparam add_49683_7.INIT1 = 16'h56aa;
    defparam add_49683_7.INJECT1_0 = "NO";
    defparam add_49683_7.INJECT1_1 = "NO";
    CCU2D add_49683_5 (.A0(n61292[3]), .B0(n12), .C0(n5), .D0(counter[3]), 
          .A1(n61292[4]), .B1(n12), .C1(n5), .D1(counter[4]), .CIN(n62584), 
          .COUT(n62585), .S0(n61278[3]), .S1(n61278[4]));
    defparam add_49683_5.INIT0 = 16'h56aa;
    defparam add_49683_5.INIT1 = 16'h56aa;
    defparam add_49683_5.INJECT1_0 = "NO";
    defparam add_49683_5.INJECT1_1 = "NO";
    LUT4 select_455_Select_2_i32_2_lut (.A(sram_output_B[2]), .B(n2022[31]), 
         .Z(n32_adj_74)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_2_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_6 (.A(\mlp_outputs[1] [2]), .B(n70809), .C(float_alu_c[2]), 
         .D(o[0]), .Z(n23216)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_6.init = 16'hc088;
    LUT4 i1_4_lut_adj_7 (.A(n32_adj_74), .B(\mlp_outputs[1] [2]), .C(n23216), 
         .D(n2022[39]), .Z(n66306)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_7.init = 16'hfefa;
    FD1P3IX o_4661__i13 (.D(n134_adj_404[13]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[13]));
    defparam o_4661__i13.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i10 (.D(\hidden_outputs[0] [10]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [10]));
    defparam temp_outputs_0__i0_i10.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i9 (.D(\hidden_outputs[0] [9]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [9]));
    defparam temp_outputs_0__i0_i9.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i8 (.D(\hidden_outputs[0] [8]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [8]));
    defparam temp_outputs_0__i0_i8.GSR = "DISABLED";
    LUT4 select_456_Select_3_i32_2_lut (.A(sram_output_B[3]), .B(n2022[31]), 
         .Z(n32_adj_75)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_3_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_8 (.A(\mlp_outputs[1] [3]), .B(n70809), .C(float_alu_c[3]), 
         .D(o[0]), .Z(n22554)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_8.init = 16'hc088;
    CCU2D add_49683_3 (.A0(n61292[1]), .B0(n12), .C0(n5), .D0(counter[1]), 
          .A1(n61292[2]), .B1(n12), .C1(n5), .D1(counter[2]), .CIN(n62583), 
          .COUT(n62584), .S0(n61278[1]), .S1(n61278[2]));
    defparam add_49683_3.INIT0 = 16'h56aa;
    defparam add_49683_3.INIT1 = 16'h55a9;
    defparam add_49683_3.INJECT1_0 = "NO";
    defparam add_49683_3.INJECT1_1 = "NO";
    FD1P3IX o_4661__i12 (.D(n134_adj_404[12]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[12]));
    defparam o_4661__i12.GSR = "DISABLED";
    FD1P3IX o_4661__i11 (.D(n134_adj_404[11]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[11]));
    defparam o_4661__i11.GSR = "DISABLED";
    FD1P3IX o_4661__i10 (.D(n134_adj_404[10]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[10]));
    defparam o_4661__i10.GSR = "DISABLED";
    CCU2D add_49683_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n61292[0]), .B1(n12), .C1(n5), .D1(counter[0]), .COUT(n62583), 
          .S1(n61278[0]));
    defparam add_49683_1.INIT0 = 16'hF000;
    defparam add_49683_1.INIT1 = 16'h55a9;
    defparam add_49683_1.INJECT1_0 = "NO";
    defparam add_49683_1.INJECT1_1 = "NO";
    FD1P3IX o_4661__i9 (.D(n134_adj_404[9]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[9]));
    defparam o_4661__i9.GSR = "DISABLED";
    FD1P3IX o_4661__i8 (.D(n134_adj_404[8]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[8]));
    defparam o_4661__i8.GSR = "DISABLED";
    FD1P3IX o_4661__i7 (.D(n134_adj_404[7]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[7]));
    defparam o_4661__i7.GSR = "DISABLED";
    FD1P3IX o_4661__i6 (.D(n134_adj_404[6]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[6]));
    defparam o_4661__i6.GSR = "DISABLED";
    FD1P3IX o_4661__i5 (.D(n134_adj_404[5]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[5]));
    defparam o_4661__i5.GSR = "DISABLED";
    FD1P3IX o_4661__i4 (.D(n134_adj_404[4]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[4]));
    defparam o_4661__i4.GSR = "DISABLED";
    FD1P3IX o_4661__i3 (.D(n134_adj_404[3]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[3]));
    defparam o_4661__i3.GSR = "DISABLED";
    FD1P3IX o_4661__i2 (.D(n134_adj_404[2]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[2]));
    defparam o_4661__i2.GSR = "DISABLED";
    FD1P3IX o_4661__i1 (.D(n134_adj_404[1]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[1]));
    defparam o_4661__i1.GSR = "DISABLED";
    LUT4 i8_2_lut (.A(numL[22]), .B(numL[24]), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    FD1P3IX counter_4663_4767__i12 (.D(n54[11]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[11]));
    defparam counter_4663_4767__i12.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i11 (.D(n54[10]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[10]));
    defparam counter_4663_4767__i11.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i10 (.D(n54[9]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[9]));
    defparam counter_4663_4767__i10.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i9 (.D(n54[8]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[8]));
    defparam counter_4663_4767__i9.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i8 (.D(n54[7]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[7]));
    defparam counter_4663_4767__i8.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i7 (.D(n54[6]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[6]));
    defparam counter_4663_4767__i7.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i6 (.D(n54[5]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[5]));
    defparam counter_4663_4767__i6.GSR = "DISABLED";
    CCU2D add_6598_12 (.A0(counter[11]), .B0(n[10]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62582), 
          .S0(n3_adj_406[11]));
    defparam add_6598_12.INIT0 = 16'h5666;
    defparam add_6598_12.INIT1 = 16'h0000;
    defparam add_6598_12.INJECT1_0 = "NO";
    defparam add_6598_12.INJECT1_1 = "NO";
    FD1P3IX counter_4663_4767__i5 (.D(n54[4]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[4]));
    defparam counter_4663_4767__i5.GSR = "DISABLED";
    FD1P3JX counter_4663_4767__i4 (.D(n54[3]), .SP(n4613), .PD(n34857), 
            .CK(clock), .Q(counter[3]));
    defparam counter_4663_4767__i4.GSR = "DISABLED";
    FD1P3JX counter_4663_4767__i3 (.D(n54[2]), .SP(n4613), .PD(n34857), 
            .CK(clock), .Q(counter[2]));
    defparam counter_4663_4767__i3.GSR = "DISABLED";
    FD1P3IX counter_4663_4767__i2 (.D(n54[1]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[1]));
    defparam counter_4663_4767__i2.GSR = "DISABLED";
    CCU2D add_6598_10 (.A0(counter[9]), .B0(n[8]), .C0(GND_net), .D0(GND_net), 
          .A1(counter[10]), .B1(n[9]), .C1(GND_net), .D1(GND_net), .CIN(n62581), 
          .COUT(n62582), .S0(n3_adj_406[9]), .S1(n3_adj_406[10]));
    defparam add_6598_10.INIT0 = 16'h5666;
    defparam add_6598_10.INIT1 = 16'h5666;
    defparam add_6598_10.INJECT1_0 = "NO";
    defparam add_6598_10.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_9 (.A(n32_adj_75), .B(n22554), .C(\mlp_outputs[1] [3]), 
         .D(n2022[39]), .Z(n66530)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_9.init = 16'hfeee;
    LUT4 i22_4_lut (.A(n31), .B(n44), .C(n40), .D(n32), .Z(n66671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 select_455_Select_4_i32_2_lut (.A(sram_output_B[4]), .B(n2022[31]), 
         .Z(n32_adj_76)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_4_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_10 (.A(\mlp_outputs[1] [4]), .B(n70809), .C(float_alu_c[4]), 
         .D(o[0]), .Z(n23174)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_10.init = 16'hc088;
    LUT4 i2_4_lut_adj_11 (.A(n23174), .B(n32_adj_76), .C(\mlp_outputs[1] [4]), 
         .D(n2022[39]), .Z(n63047)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_11.init = 16'hfeee;
    LUT4 i112_3_lut_4_lut (.A(h[0]), .B(n70847), .C(n2448[31]), .D(\hidden_outputs[0] [31]), 
         .Z(n1586)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C))) */ ;
    defparam i112_3_lut_4_lut.init = 16'hef01;
    CCU2D add_6598_8 (.A0(counter[7]), .B0(n[6]), .C0(GND_net), .D0(GND_net), 
          .A1(counter[8]), .B1(n[7]), .C1(GND_net), .D1(GND_net), .CIN(n62580), 
          .COUT(n62581), .S0(n3_adj_406[7]), .S1(n3_adj_406[8]));
    defparam add_6598_8.INIT0 = 16'h5666;
    defparam add_6598_8.INIT1 = 16'h5666;
    defparam add_6598_8.INJECT1_0 = "NO";
    defparam add_6598_8.INJECT1_1 = "NO";
    CCU2D add_6598_6 (.A0(counter[5]), .B0(n[4]), .C0(GND_net), .D0(GND_net), 
          .A1(counter[6]), .B1(n[5]), .C1(GND_net), .D1(GND_net), .CIN(n62579), 
          .COUT(n62580), .S0(n3_adj_406[5]), .S1(n3_adj_406[6]));
    defparam add_6598_6.INIT0 = 16'h5666;
    defparam add_6598_6.INIT1 = 16'h5666;
    defparam add_6598_6.INJECT1_0 = "NO";
    defparam add_6598_6.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_12 (.A(\hidden_outputs[4] [0]), .B(n22568), .C(float_alu_c[0]), 
         .D(n70783), .Z(n22745)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_12.init = 16'hc088;
    CCU2D add_6598_4 (.A0(counter[3]), .B0(n[2]), .C0(GND_net), .D0(GND_net), 
          .A1(counter[4]), .B1(n[3]), .C1(GND_net), .D1(GND_net), .CIN(n62578), 
          .COUT(n62579), .S0(n3_adj_406[3]), .S1(n3_adj_406[4]));
    defparam add_6598_4.INIT0 = 16'h5666;
    defparam add_6598_4.INIT1 = 16'h5666;
    defparam add_6598_4.INJECT1_0 = "NO";
    defparam add_6598_4.INJECT1_1 = "NO";
    CCU2D add_6598_2 (.A0(counter[1]), .B0(n[0]), .C0(GND_net), .D0(GND_net), 
          .A1(counter[2]), .B1(n[1]), .C1(GND_net), .D1(GND_net), .COUT(n62578), 
          .S1(n3_adj_406[2]));
    defparam add_6598_2.INIT0 = 16'h7000;
    defparam add_6598_2.INIT1 = 16'h5666;
    defparam add_6598_2.INJECT1_0 = "NO";
    defparam add_6598_2.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_13 (.A(n10_adj_77), .B(n22745), .C(\hidden_outputs[4] [0]), 
         .D(n2022[17]), .Z(n66466)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_13.init = 16'hfeee;
    CCU2D add_49682_12 (.A0(n3[10]), .B0(n70712), .C0(h[10]), .D0(n7729[9]), 
          .A1(n3[11]), .B1(n70712), .C1(h[11]), .D1(n7729[10]), .CIN(n62575), 
          .S0(n61264[10]), .S1(n61264[11]));
    defparam add_49682_12.INIT0 = 16'h596a;
    defparam add_49682_12.INIT1 = 16'h596a;
    defparam add_49682_12.INJECT1_0 = "NO";
    defparam add_49682_12.INJECT1_1 = "NO";
    LUT4 select_456_Select_5_i32_2_lut (.A(sram_output_B[5]), .B(n2022[31]), 
         .Z(n32_adj_80)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_5_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_14 (.A(\mlp_outputs[1] [5]), .B(n70809), .C(float_alu_c[5]), 
         .D(o[0]), .Z(n22742)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_14.init = 16'hc088;
    LUT4 i1_4_lut_adj_15 (.A(n32_adj_80), .B(n22742), .C(\mlp_outputs[1] [5]), 
         .D(n2022[39]), .Z(n66468)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_15.init = 16'hfeee;
    FD1P3AX temp_outputs_1__i0_i24 (.D(\hidden_outputs[1] [24]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [24]));
    defparam temp_outputs_1__i0_i24.GSR = "DISABLED";
    LUT4 i4_4_lut (.A(numL[6]), .B(numL[25]), .C(numL[16]), .D(numL[3]), 
         .Z(n10_adj_81)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut.init = 16'hfffe;
    CCU2D add_49682_10 (.A0(n3[8]), .B0(n70712), .C0(h[8]), .D0(n7729[7]), 
          .A1(n3[9]), .B1(n70712), .C1(h[9]), .D1(n7729[8]), .CIN(n62574), 
          .COUT(n62575), .S0(n61264[8]), .S1(n61264[9]));
    defparam add_49682_10.INIT0 = 16'h596a;
    defparam add_49682_10.INIT1 = 16'h596a;
    defparam add_49682_10.INJECT1_0 = "NO";
    defparam add_49682_10.INJECT1_1 = "NO";
    LUT4 select_455_Select_6_i32_2_lut (.A(sram_output_B[6]), .B(n2022[31]), 
         .Z(n32_adj_84)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_6_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_16 (.A(\mlp_outputs[1] [6]), .B(n70809), .C(float_alu_c[6]), 
         .D(o[0]), .Z(n23240)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_16.init = 16'hc088;
    LUT4 i1_4_lut_adj_17 (.A(n32_adj_84), .B(\mlp_outputs[1] [6]), .C(n23240), 
         .D(n2022[39]), .Z(n66292)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_17.init = 16'hfefa;
    CCU2D add_49682_8 (.A0(n3[6]), .B0(n70712), .C0(h[6]), .D0(n7729[5]), 
          .A1(n3[7]), .B1(n70712), .C1(h[7]), .D1(n7729[6]), .CIN(n62573), 
          .COUT(n62574), .S0(n61264[6]), .S1(n61264[7]));
    defparam add_49682_8.INIT0 = 16'h596a;
    defparam add_49682_8.INIT1 = 16'h596a;
    defparam add_49682_8.INJECT1_0 = "NO";
    defparam add_49682_8.INJECT1_1 = "NO";
    LUT4 select_460_Select_0_i94_2_lut (.A(n2022[22]), .B(n2022[24]), .Z(n17400)) /* synthesis lut_function=(A+(B)) */ ;
    defparam select_460_Select_0_i94_2_lut.init = 16'heeee;
    CCU2D add_49682_6 (.A0(n3[4]), .B0(n70712), .C0(h[4]), .D0(n7729[3]), 
          .A1(n3[5]), .B1(n70712), .C1(h[5]), .D1(n7729[4]), .CIN(n62572), 
          .COUT(n62573), .S0(n61264[4]), .S1(n61264[5]));
    defparam add_49682_6.INIT0 = 16'h596a;
    defparam add_49682_6.INIT1 = 16'h596a;
    defparam add_49682_6.INJECT1_0 = "NO";
    defparam add_49682_6.INJECT1_1 = "NO";
    CCU2D add_49682_4 (.A0(n3[2]), .B0(n70712), .C0(h[2]), .D0(n7729[1]), 
          .A1(n3[3]), .B1(n70712), .C1(h[3]), .D1(n7729[2]), .CIN(n62571), 
          .COUT(n62572), .S0(n61264[2]), .S1(n61264[3]));
    defparam add_49682_4.INIT0 = 16'h596a;
    defparam add_49682_4.INIT1 = 16'h596a;
    defparam add_49682_4.INJECT1_0 = "NO";
    defparam add_49682_4.INJECT1_1 = "NO";
    CCU2D add_49682_2 (.A0(n3[0]), .B0(h[0]), .C0(GND_net), .D0(GND_net), 
          .A1(n3[1]), .B1(i[0]), .C1(n70712), .D1(h[1]), .COUT(n62571), 
          .S1(n61264[1]));
    defparam add_49682_2.INIT0 = 16'h7000;
    defparam add_49682_2.INIT1 = 16'h59a6;
    defparam add_49682_2.INJECT1_0 = "NO";
    defparam add_49682_2.INJECT1_1 = "NO";
    LUT4 i55072_3_lut_4_lut (.A(h[0]), .B(n70847), .C(n40754), .D(n2022[9]), 
         .Z(n23658)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i55072_3_lut_4_lut.init = 16'h10f0;
    LUT4 i7063_2_lut (.A(i[0]), .B(i[1]), .Z(n17802)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7063_2_lut.init = 16'heeee;
    LUT4 mux_75_Mux_0_i7_4_lut (.A(n67260), .B(\temp_outputs[4] [0]), .C(i[2]), 
         .D(n17802), .Z(n1028[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_0_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i1_3_lut (.A(n1028[0]), .B(n1027[0]), .C(n70712), .Z(n1061[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i1_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_18 (.A(f[0]), .B(n2448[0]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_89)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_18.init = 16'heca0;
    LUT4 select_460_Select_0_i16_2_lut (.A(e[0]), .B(n2022[15]), .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_0_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_19 (.A(n18717), .B(n8_adj_89), .C(n1061[0]), .D(n2022[13]), 
         .Z(n10_adj_90)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_19.init = 16'hfeee;
    CCU2D add_49681_13 (.A0(n61264[11]), .B0(n12), .C0(n5), .D0(counter[11]), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62569), 
          .S0(n61250[11]));
    defparam add_49681_13.INIT0 = 16'h56aa;
    defparam add_49681_13.INIT1 = 16'h0000;
    defparam add_49681_13.INJECT1_0 = "NO";
    defparam add_49681_13.INJECT1_1 = "NO";
    CCU2D add_49681_11 (.A0(n61264[9]), .B0(n12), .C0(n5), .D0(counter[9]), 
          .A1(n61264[10]), .B1(n12), .C1(n5), .D1(counter[10]), .CIN(n62568), 
          .COUT(n62569), .S0(n61250[9]), .S1(n61250[10]));
    defparam add_49681_11.INIT0 = 16'h56aa;
    defparam add_49681_11.INIT1 = 16'h56aa;
    defparam add_49681_11.INJECT1_0 = "NO";
    defparam add_49681_11.INJECT1_1 = "NO";
    LUT4 mux_220_Mux_0_i7_4_lut (.A(n67254), .B(\hidden_outputs[4] [0]), 
         .C(n[2]), .D(n70842), .Z(n3742[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_0_i7_4_lut.init = 16'h0aca;
    CCU2D add_49681_9 (.A0(n61264[7]), .B0(n12), .C0(n5), .D0(counter[7]), 
          .A1(n61264[8]), .B1(n12), .C1(n5), .D1(counter[8]), .CIN(n62567), 
          .COUT(n62568), .S0(n61250[7]), .S1(n61250[8]));
    defparam add_49681_9.INIT0 = 16'h56aa;
    defparam add_49681_9.INIT1 = 16'h56aa;
    defparam add_49681_9.INJECT1_0 = "NO";
    defparam add_49681_9.INJECT1_1 = "NO";
    CCU2D add_49681_7 (.A0(n61264[5]), .B0(n12), .C0(n5), .D0(counter[5]), 
          .A1(n61264[6]), .B1(n12), .C1(n5), .D1(counter[6]), .CIN(n62566), 
          .COUT(n62567), .S0(n61250[5]), .S1(n61250[6]));
    defparam add_49681_7.INIT0 = 16'h56aa;
    defparam add_49681_7.INIT1 = 16'h56aa;
    defparam add_49681_7.INJECT1_0 = "NO";
    defparam add_49681_7.INJECT1_1 = "NO";
    LUT4 i5_4_lut (.A(n3742[0]), .B(n10_adj_90), .C(n16), .D(n2022[35]), 
         .Z(n63022)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    CCU2D add_49681_5 (.A0(n61264[3]), .B0(n12), .C0(n5), .D0(counter[3]), 
          .A1(n61264[4]), .B1(n12), .C1(n5), .D1(counter[4]), .CIN(n62565), 
          .COUT(n62566), .S0(n61250[3]), .S1(n61250[4]));
    defparam add_49681_5.INIT0 = 16'h56aa;
    defparam add_49681_5.INIT1 = 16'h56aa;
    defparam add_49681_5.INJECT1_0 = "NO";
    defparam add_49681_5.INJECT1_1 = "NO";
    CCU2D add_49681_3 (.A0(n61264[1]), .B0(n12), .C0(n5), .D0(counter[1]), 
          .A1(n61264[2]), .B1(n12), .C1(n5), .D1(counter[2]), .CIN(n62564), 
          .COUT(n62565), .S0(n61250[1]), .S1(n61250[2]));
    defparam add_49681_3.INIT0 = 16'h56aa;
    defparam add_49681_3.INIT1 = 16'h55a9;
    defparam add_49681_3.INJECT1_0 = "NO";
    defparam add_49681_3.INJECT1_1 = "NO";
    CCU2D add_49681_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n61264[0]), .B1(n12), .C1(n5), .D1(counter[0]), .COUT(n62564), 
          .S1(n61250[0]));
    defparam add_49681_1.INIT0 = 16'hF000;
    defparam add_49681_1.INIT1 = 16'h55a9;
    defparam add_49681_1.INJECT1_0 = "NO";
    defparam add_49681_1.INJECT1_1 = "NO";
    FD1P3AX temp_outputs_1__i0_i26 (.D(\hidden_outputs[1] [26]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[1] [26]));
    defparam temp_outputs_1__i0_i26.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i7 (.D(\hidden_outputs[0] [7]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [7]));
    defparam temp_outputs_0__i0_i7.GSR = "DISABLED";
    LUT4 i111_3_lut_4_lut (.A(h[0]), .B(n70847), .C(n2448[31]), .D(\hidden_outputs[1] [31]), 
         .Z(n1585)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (D)) */ ;
    defparam i111_3_lut_4_lut.init = 16'hdf02;
    LUT4 i55053_3_lut_4_lut (.A(h[0]), .B(n70847), .C(n40754), .D(n2022[9]), 
         .Z(n23659)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;
    defparam i55053_3_lut_4_lut.init = 16'h20f0;
    LUT4 i1_4_lut_adj_20 (.A(\hidden_outputs[3] [0]), .B(n22568), .C(float_alu_c[0]), 
         .D(n70785), .Z(n23363)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_20.init = 16'hc088;
    LUT4 i1_4_lut_adj_21 (.A(n10_adj_77), .B(\hidden_outputs[3] [0]), .C(n23363), 
         .D(n2022[17]), .Z(n66386)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_21.init = 16'hfefa;
    PFUMX i54343 (.BLUT(n67252), .ALUT(n67253), .C0(n[1]), .Z(n67254));
    CCU2D add_3865_13 (.A0(o[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62549), 
          .S0(n11102[11]));
    defparam add_3865_13.INIT0 = 16'hfaaa;
    defparam add_3865_13.INIT1 = 16'h0000;
    defparam add_3865_13.INJECT1_0 = "NO";
    defparam add_3865_13.INJECT1_1 = "NO";
    LUT4 select_456_Select_7_i32_2_lut (.A(sram_output_B[7]), .B(n2022[31]), 
         .Z(n32_adj_91)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_7_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_22 (.A(\mlp_outputs[1] [7]), .B(n70809), .C(float_alu_c[7]), 
         .D(o[0]), .Z(n23237)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_22.init = 16'hc088;
    LUT4 i2_4_lut_adj_23 (.A(n23237), .B(n32_adj_91), .C(\mlp_outputs[1] [7]), 
         .D(n2022[39]), .Z(n63058)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_23.init = 16'hfeee;
    CCU2D add_3865_11 (.A0(o[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62548), 
          .COUT(n62549), .S0(n11102[9]), .S1(n11102[10]));
    defparam add_3865_11.INIT0 = 16'hfaaa;
    defparam add_3865_11.INIT1 = 16'hfaaa;
    defparam add_3865_11.INJECT1_0 = "NO";
    defparam add_3865_11.INJECT1_1 = "NO";
    CCU2D add_3865_9 (.A0(o[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62547), 
          .COUT(n62548), .S0(n11102[7]), .S1(n11102[8]));
    defparam add_3865_9.INIT0 = 16'hfaaa;
    defparam add_3865_9.INIT1 = 16'hfaaa;
    defparam add_3865_9.INJECT1_0 = "NO";
    defparam add_3865_9.INJECT1_1 = "NO";
    CCU2D add_3865_7 (.A0(o[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62546), 
          .COUT(n62547), .S0(n11102[5]), .S1(n11102[6]));
    defparam add_3865_7.INIT0 = 16'hfaaa;
    defparam add_3865_7.INIT1 = 16'hfaaa;
    defparam add_3865_7.INJECT1_0 = "NO";
    defparam add_3865_7.INJECT1_1 = "NO";
    CCU2D add_3865_5 (.A0(o[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62545), 
          .COUT(n62546), .S0(n11102[3]), .S1(n11102[4]));
    defparam add_3865_5.INIT0 = 16'h0555;
    defparam add_3865_5.INIT1 = 16'h0555;
    defparam add_3865_5.INJECT1_0 = "NO";
    defparam add_3865_5.INJECT1_1 = "NO";
    LUT4 select_455_Select_8_i32_2_lut (.A(sram_output_B[8]), .B(n2022[31]), 
         .Z(n32_adj_92)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_8_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_24 (.A(\mlp_outputs[1] [8]), .B(n70809), .C(float_alu_c[8]), 
         .D(o[0]), .Z(n23183)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_24.init = 16'hc088;
    LUT4 i1_4_lut_adj_25 (.A(n32_adj_92), .B(\mlp_outputs[1] [8]), .C(n23183), 
         .D(n2022[39]), .Z(n66474)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_25.init = 16'hfefa;
    CCU2D add_3865_3 (.A0(o[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62544), 
          .COUT(n62545), .S0(n11102[1]), .S1(n11102[2]));
    defparam add_3865_3.INIT0 = 16'h0555;
    defparam add_3865_3.INIT1 = 16'hfaaa;
    defparam add_3865_3.INJECT1_0 = "NO";
    defparam add_3865_3.INJECT1_1 = "NO";
    CCU2D add_3865_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(o[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62544), 
          .S1(n11102[0]));
    defparam add_3865_1.INIT0 = 16'hF000;
    defparam add_3865_1.INIT1 = 16'h0555;
    defparam add_3865_1.INJECT1_0 = "NO";
    defparam add_3865_1.INJECT1_1 = "NO";
    LUT4 i54630_3_lut (.A(\hidden_outputs[2] [31]), .B(\hidden_outputs[3] [31]), 
         .C(n[0]), .Z(n67541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54630_3_lut.init = 16'hcaca;
    LUT4 i54629_3_lut (.A(\hidden_outputs[0] [31]), .B(\hidden_outputs[1] [31]), 
         .C(n[0]), .Z(n67540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54629_3_lut.init = 16'hcaca;
    LUT4 i54627_3_lut (.A(\hidden_outputs[2] [30]), .B(\hidden_outputs[3] [30]), 
         .C(n[0]), .Z(n67538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54627_3_lut.init = 16'hcaca;
    LUT4 i54626_3_lut (.A(\hidden_outputs[0] [30]), .B(\hidden_outputs[1] [30]), 
         .C(n[0]), .Z(n67537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54626_3_lut.init = 16'hcaca;
    LUT4 i54624_3_lut (.A(\hidden_outputs[2] [29]), .B(\hidden_outputs[3] [29]), 
         .C(n[0]), .Z(n67535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54624_3_lut.init = 16'hcaca;
    LUT4 i54623_3_lut (.A(\hidden_outputs[0] [29]), .B(\hidden_outputs[1] [29]), 
         .C(n[0]), .Z(n67534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54623_3_lut.init = 16'hcaca;
    LUT4 select_455_Select_9_i32_2_lut (.A(sram_output_B[9]), .B(n2022[31]), 
         .Z(n32_adj_93)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_9_i32_2_lut.init = 16'h8888;
    LUT4 i55048_3_lut_4_lut (.A(h[0]), .B(n70845), .C(n40754), .D(n2022[9]), 
         .Z(n23660)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;
    defparam i55048_3_lut_4_lut.init = 16'h40f0;
    LUT4 i54621_3_lut (.A(\hidden_outputs[2] [28]), .B(\hidden_outputs[3] [28]), 
         .C(n[0]), .Z(n67532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54621_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_26 (.A(\mlp_outputs[1] [9]), .B(n70809), .C(float_alu_c[9]), 
         .D(o[0]), .Z(n23483)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_26.init = 16'hc088;
    LUT4 i1_4_lut_adj_27 (.A(n32_adj_93), .B(\mlp_outputs[1] [9]), .C(n23483), 
         .D(n2022[39]), .Z(n66348)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_27.init = 16'hfefa;
    LUT4 i110_3_lut_4_lut (.A(h[0]), .B(n70845), .C(n2448[31]), .D(\hidden_outputs[2] [31]), 
         .Z(n1584)) /* synthesis lut_function=(A (D)+!A !(B (C)+!B !(D))) */ ;
    defparam i110_3_lut_4_lut.init = 16'hbf04;
    LUT4 i54620_3_lut (.A(\hidden_outputs[0] [28]), .B(\hidden_outputs[1] [28]), 
         .C(n[0]), .Z(n67531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54620_3_lut.init = 16'hcaca;
    LUT4 i54618_3_lut (.A(\hidden_outputs[2] [27]), .B(\hidden_outputs[3] [27]), 
         .C(n[0]), .Z(n67529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54618_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_761_4_lut (.A(numL[18]), .B(n10_adj_81), .C(numL[7]), 
         .D(n66671), .Z(n70731)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_761_4_lut.init = 16'hfffe;
    LUT4 i54617_3_lut (.A(\hidden_outputs[0] [27]), .B(\hidden_outputs[1] [27]), 
         .C(n[0]), .Z(n67528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54617_3_lut.init = 16'hcaca;
    LUT4 i5_3_lut_rep_816 (.A(numL[18]), .B(n10_adj_81), .C(numL[7]), 
         .Z(n70786)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut_rep_816.init = 16'hfefe;
    LUT4 i1_2_lut_adj_28 (.A(n23104), .B(n2448[24]), .Z(n23327)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_28.init = 16'h8888;
    LUT4 i2_4_lut_adj_29 (.A(n23327), .B(n23330), .C(weight[24]), .D(n70860), 
         .Z(n63111)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_29.init = 16'hfeee;
    LUT4 i109_3_lut_4_lut (.A(h[0]), .B(n70845), .C(n2448[31]), .D(\hidden_outputs[3] [31]), 
         .Z(n1583)) /* synthesis lut_function=(!(A (B (C)+!B !(D))+!A !(D))) */ ;
    defparam i109_3_lut_4_lut.init = 16'h7f08;
    LUT4 i54615_3_lut (.A(\hidden_outputs[2] [26]), .B(\hidden_outputs[3] [26]), 
         .C(n[0]), .Z(n67526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54615_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_30 (.A(mlp_mode), .B(mlp_ready), .Z(n23661)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_30.init = 16'h4444;
    LUT4 i55102_3_lut_4_lut (.A(h[0]), .B(n70845), .C(n40754), .D(n2022[9]), 
         .Z(n23663)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i55102_3_lut_4_lut.init = 16'h80f0;
    LUT4 i108_3_lut_4_lut (.A(h[2]), .B(n70861), .C(n2448[31]), .D(\hidden_outputs[4] [31]), 
         .Z(n1582)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (D)) */ ;
    defparam i108_3_lut_4_lut.init = 16'hdf02;
    LUT4 i55100_3_lut_4_lut (.A(h[2]), .B(n70861), .C(n40754), .D(n2022[9]), 
         .Z(n23665)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;
    defparam i55100_3_lut_4_lut.init = 16'h20f0;
    FD1P3DX float_alu_mode_i0_i1 (.D(n23977), .SP(n27939), .CK(clock), 
            .CD(SDA_c), .Q(\float_alu_mode[1] ));
    defparam float_alu_mode_i0_i1.GSR = "DISABLED";
    LUT4 i54614_3_lut (.A(\hidden_outputs[0] [26]), .B(\hidden_outputs[1] [26]), 
         .C(n[0]), .Z(n67525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54614_3_lut.init = 16'hcaca;
    LUT4 i54612_3_lut (.A(\hidden_outputs[2] [25]), .B(\hidden_outputs[3] [25]), 
         .C(n[0]), .Z(n67523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54612_3_lut.init = 16'hcaca;
    LUT4 i54611_3_lut (.A(\hidden_outputs[0] [25]), .B(\hidden_outputs[1] [25]), 
         .C(n[0]), .Z(n67522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54611_3_lut.init = 16'hcaca;
    LUT4 i54609_3_lut (.A(\hidden_outputs[2] [24]), .B(\hidden_outputs[3] [24]), 
         .C(n[0]), .Z(n67520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54609_3_lut.init = 16'hcaca;
    LUT4 i54608_3_lut (.A(\hidden_outputs[0] [24]), .B(\hidden_outputs[1] [24]), 
         .C(n[0]), .Z(n67519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54608_3_lut.init = 16'hcaca;
    LUT4 i54606_3_lut (.A(\hidden_outputs[2] [23]), .B(\hidden_outputs[3] [23]), 
         .C(n[0]), .Z(n67517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54606_3_lut.init = 16'hcaca;
    LUT4 i54605_3_lut (.A(\hidden_outputs[0] [23]), .B(\hidden_outputs[1] [23]), 
         .C(n[0]), .Z(n67516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54605_3_lut.init = 16'hcaca;
    LUT4 select_455_Select_10_i32_2_lut (.A(sram_output_B[10]), .B(n2022[31]), 
         .Z(n32_adj_94)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_10_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_31 (.A(\mlp_outputs[1] [10]), .B(n70809), .C(float_alu_c[10]), 
         .D(o[0]), .Z(n23297)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_31.init = 16'hc088;
    LUT4 i1_2_lut_adj_32 (.A(n23104), .B(n2448[26]), .Z(n81)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_32.init = 16'h8888;
    LUT4 i1_4_lut_adj_33 (.A(n32_adj_94), .B(\mlp_outputs[1] [10]), .C(n23297), 
         .D(n2022[39]), .Z(n66526)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_33.init = 16'hfefa;
    LUT4 i2_4_lut_adj_34 (.A(n81), .B(n23339), .C(weight[26]), .D(n70860), 
         .Z(n63112)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_34.init = 16'hfeee;
    LUT4 i54603_3_lut (.A(\hidden_outputs[2] [22]), .B(\hidden_outputs[3] [22]), 
         .C(n[0]), .Z(n67514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54603_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_35 (.A(\hidden_outputs[2] [0]), .B(n22568), .C(float_alu_c[0]), 
         .D(n70787), .Z(n22937)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_35.init = 16'hc088;
    LUT4 i54602_3_lut (.A(\hidden_outputs[0] [22]), .B(\hidden_outputs[1] [22]), 
         .C(n[0]), .Z(n67513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54602_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_36 (.A(n10_adj_77), .B(n22937), .C(\hidden_outputs[2] [0]), 
         .D(n2022[17]), .Z(n66300)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_36.init = 16'hfeee;
    LUT4 i54600_3_lut (.A(\hidden_outputs[2] [21]), .B(\hidden_outputs[3] [21]), 
         .C(n[0]), .Z(n67511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54600_3_lut.init = 16'hcaca;
    LUT4 select_455_Select_11_i32_2_lut (.A(sram_output_B[11]), .B(n2022[31]), 
         .Z(n32_adj_95)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_11_i32_2_lut.init = 16'h8888;
    LUT4 i54599_3_lut (.A(\hidden_outputs[0] [21]), .B(\hidden_outputs[1] [21]), 
         .C(n[0]), .Z(n67510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54599_3_lut.init = 16'hcaca;
    LUT4 i54597_3_lut (.A(\hidden_outputs[2] [20]), .B(\hidden_outputs[3] [20]), 
         .C(n[0]), .Z(n67508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54597_3_lut.init = 16'hcaca;
    LUT4 i54596_3_lut (.A(\hidden_outputs[0] [20]), .B(\hidden_outputs[1] [20]), 
         .C(n[0]), .Z(n67507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54596_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_37 (.A(\mlp_outputs[1] [11]), .B(n70809), .C(float_alu_c[11]), 
         .D(o[0]), .Z(n23186)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_37.init = 16'hc088;
    LUT4 i54594_3_lut (.A(\hidden_outputs[2] [19]), .B(\hidden_outputs[3] [19]), 
         .C(n[0]), .Z(n67505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54594_3_lut.init = 16'hcaca;
    LUT4 i54593_3_lut (.A(\hidden_outputs[0] [19]), .B(\hidden_outputs[1] [19]), 
         .C(n[0]), .Z(n67504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54593_3_lut.init = 16'hcaca;
    LUT4 i54591_3_lut (.A(\hidden_outputs[2] [18]), .B(\hidden_outputs[3] [18]), 
         .C(n[0]), .Z(n67502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54591_3_lut.init = 16'hcaca;
    LUT4 i54590_3_lut (.A(\hidden_outputs[0] [18]), .B(\hidden_outputs[1] [18]), 
         .C(n[0]), .Z(n67501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54590_3_lut.init = 16'hcaca;
    LUT4 i54588_3_lut (.A(\hidden_outputs[2] [17]), .B(\hidden_outputs[3] [17]), 
         .C(n[0]), .Z(n67499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54588_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_38 (.A(n32_adj_95), .B(\mlp_outputs[1] [11]), .C(n23186), 
         .D(n2022[39]), .Z(n66400)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_38.init = 16'hfefa;
    LUT4 select_455_Select_12_i32_2_lut (.A(sram_output_B[12]), .B(n2022[31]), 
         .Z(n32_adj_96)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_12_i32_2_lut.init = 16'h8888;
    LUT4 i54587_3_lut (.A(\hidden_outputs[0] [17]), .B(\hidden_outputs[1] [17]), 
         .C(n[0]), .Z(n67498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54587_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_39 (.A(\mlp_outputs[1] [12]), .B(n70809), .C(float_alu_c[12]), 
         .D(o[0]), .Z(n23321)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_39.init = 16'hc088;
    LUT4 i54585_3_lut (.A(\hidden_outputs[2] [16]), .B(\hidden_outputs[3] [16]), 
         .C(n[0]), .Z(n67496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54585_3_lut.init = 16'hcaca;
    LUT4 i54584_3_lut (.A(\hidden_outputs[0] [16]), .B(\hidden_outputs[1] [16]), 
         .C(n[0]), .Z(n67495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54584_3_lut.init = 16'hcaca;
    LUT4 i54582_3_lut (.A(\hidden_outputs[2] [15]), .B(\hidden_outputs[3] [15]), 
         .C(n[0]), .Z(n67493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54582_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_40 (.A(n32_adj_96), .B(\mlp_outputs[1] [12]), .C(n23321), 
         .D(n2022[39]), .Z(n66390)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_40.init = 16'hfefa;
    LUT4 select_455_Select_13_i32_2_lut (.A(sram_output_B[13]), .B(n2022[31]), 
         .Z(n32_adj_97)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_13_i32_2_lut.init = 16'h8888;
    LUT4 i54581_3_lut (.A(\hidden_outputs[0] [15]), .B(\hidden_outputs[1] [15]), 
         .C(n[0]), .Z(n67492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54581_3_lut.init = 16'hcaca;
    LUT4 i54579_3_lut (.A(\hidden_outputs[2] [14]), .B(\hidden_outputs[3] [14]), 
         .C(n[0]), .Z(n67490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54579_3_lut.init = 16'hcaca;
    LUT4 i54578_3_lut (.A(\hidden_outputs[0] [14]), .B(\hidden_outputs[1] [14]), 
         .C(n[0]), .Z(n67489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54578_3_lut.init = 16'hcaca;
    LUT4 i54576_3_lut (.A(\hidden_outputs[2] [13]), .B(\hidden_outputs[3] [13]), 
         .C(n[0]), .Z(n67487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54576_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_41 (.A(\mlp_outputs[1] [13]), .B(n70809), .C(float_alu_c[13]), 
         .D(o[0]), .Z(n22772)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_41.init = 16'hc088;
    LUT4 i54575_3_lut (.A(\hidden_outputs[0] [13]), .B(\hidden_outputs[1] [13]), 
         .C(n[0]), .Z(n67486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54575_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_42 (.A(n32_adj_97), .B(n22772), .C(\mlp_outputs[1] [13]), 
         .D(n2022[39]), .Z(n66460)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_42.init = 16'hfeee;
    LUT4 select_455_Select_14_i32_2_lut (.A(sram_output_B[14]), .B(n2022[31]), 
         .Z(n32_adj_98)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_14_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_43 (.A(\mlp_outputs[1] [14]), .B(n70809), .C(float_alu_c[14]), 
         .D(o[0]), .Z(n22775)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_43.init = 16'hc088;
    LUT4 i54573_3_lut (.A(\hidden_outputs[2] [12]), .B(\hidden_outputs[3] [12]), 
         .C(n[0]), .Z(n67484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54573_3_lut.init = 16'hcaca;
    LUT4 i54572_3_lut (.A(\hidden_outputs[0] [12]), .B(\hidden_outputs[1] [12]), 
         .C(n[0]), .Z(n67483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54572_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_44 (.A(n32_adj_98), .B(n22775), .C(\mlp_outputs[1] [14]), 
         .D(n2022[39]), .Z(n66458)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_44.init = 16'hfeee;
    LUT4 select_455_Select_15_i32_2_lut (.A(sram_output_B[15]), .B(n2022[31]), 
         .Z(n32_adj_99)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_15_i32_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_766_4_lut (.A(n70857), .B(n70812), .C(n128), .D(n22276), 
         .Z(n70736)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_766_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_45 (.A(\mlp_outputs[1] [15]), .B(n70809), .C(float_alu_c[15]), 
         .D(o[0]), .Z(n23516)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_45.init = 16'hc088;
    LUT4 i2_4_lut_adj_46 (.A(n23516), .B(n32_adj_99), .C(\mlp_outputs[1] [15]), 
         .D(n2022[39]), .Z(n63246)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_46.init = 16'hfeee;
    LUT4 select_455_Select_16_i32_2_lut (.A(sram_output_B[16]), .B(n2022[31]), 
         .Z(n32_adj_100)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_16_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_47 (.A(\mlp_outputs[1] [16]), .B(n70809), .C(float_alu_c[16]), 
         .D(o[0]), .Z(n23513)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_47.init = 16'hc088;
    LUT4 i1_4_lut_adj_48 (.A(n32_adj_100), .B(\mlp_outputs[1] [16]), .C(n23513), 
         .D(n2022[39]), .Z(n66334)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_48.init = 16'hfefa;
    LUT4 select_455_Select_17_i32_2_lut (.A(sram_output_B[17]), .B(n2022[31]), 
         .Z(n32_adj_101)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_17_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_49 (.A(\mlp_outputs[1] [17]), .B(n70809), .C(float_alu_c[17]), 
         .D(o[0]), .Z(n22799)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_49.init = 16'hc088;
    LUT4 i1_4_lut_adj_50 (.A(n32_adj_101), .B(n22799), .C(\mlp_outputs[1] [17]), 
         .D(n2022[39]), .Z(n66456)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_50.init = 16'hfeee;
    LUT4 select_455_Select_18_i32_2_lut (.A(sram_output_B[18]), .B(n2022[31]), 
         .Z(n32_adj_102)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_18_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_51 (.A(\mlp_outputs[1] [18]), .B(n70809), .C(float_alu_c[18]), 
         .D(o[0]), .Z(n23507)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_51.init = 16'hc088;
    LUT4 i1_4_lut_adj_52 (.A(n32_adj_102), .B(\mlp_outputs[1] [18]), .C(n23507), 
         .D(n2022[39]), .Z(n66338)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_52.init = 16'hfefa;
    LUT4 select_455_Select_19_i32_2_lut (.A(sram_output_B[19]), .B(n2022[31]), 
         .Z(n32_adj_103)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_19_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_53 (.A(\mlp_outputs[1] [19]), .B(n70809), .C(float_alu_c[19]), 
         .D(o[0]), .Z(n23510)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_53.init = 16'hc088;
    LUT4 i54570_3_lut (.A(\hidden_outputs[2] [11]), .B(\hidden_outputs[3] [11]), 
         .C(n[0]), .Z(n67481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54570_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_54 (.A(n32_adj_103), .B(\mlp_outputs[1] [19]), .C(n23510), 
         .D(n2022[39]), .Z(n66336)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_54.init = 16'hfefa;
    LUT4 i54569_3_lut (.A(\hidden_outputs[0] [11]), .B(\hidden_outputs[1] [11]), 
         .C(n[0]), .Z(n67480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54569_3_lut.init = 16'hcaca;
    LUT4 i54567_3_lut (.A(\hidden_outputs[2] [10]), .B(\hidden_outputs[3] [10]), 
         .C(n[0]), .Z(n67478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54567_3_lut.init = 16'hcaca;
    LUT4 i54566_3_lut (.A(\hidden_outputs[0] [10]), .B(\hidden_outputs[1] [10]), 
         .C(n[0]), .Z(n67477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54566_3_lut.init = 16'hcaca;
    LUT4 i49862_2_lut (.A(n2664), .B(numL[0]), .Z(n134_adj_407[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49862_2_lut.init = 16'h6666;
    LUT4 i54564_3_lut (.A(\hidden_outputs[2] [9]), .B(\hidden_outputs[3] [9]), 
         .C(n[0]), .Z(n67475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54564_3_lut.init = 16'hcaca;
    LUT4 i54563_3_lut (.A(\hidden_outputs[0] [9]), .B(\hidden_outputs[1] [9]), 
         .C(n[0]), .Z(n67474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54563_3_lut.init = 16'hcaca;
    LUT4 select_455_Select_20_i32_2_lut (.A(sram_output_B[20]), .B(n2022[31]), 
         .Z(n32_adj_105)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_20_i32_2_lut.init = 16'h8888;
    LUT4 i54561_3_lut (.A(\hidden_outputs[2] [8]), .B(\hidden_outputs[3] [8]), 
         .C(n[0]), .Z(n67472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54561_3_lut.init = 16'hcaca;
    LUT4 i54560_3_lut (.A(\hidden_outputs[0] [8]), .B(\hidden_outputs[1] [8]), 
         .C(n[0]), .Z(n67471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54560_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_55 (.A(\mlp_outputs[1] [20]), .B(n70809), .C(float_alu_c[20]), 
         .D(o[0]), .Z(n22548)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_55.init = 16'hc088;
    LUT4 i1_4_lut_adj_56 (.A(n32_adj_105), .B(n22548), .C(\mlp_outputs[1] [20]), 
         .D(n2022[39]), .Z(n66322)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_56.init = 16'hfeee;
    LUT4 i54558_3_lut (.A(\hidden_outputs[2] [7]), .B(\hidden_outputs[3] [7]), 
         .C(n[0]), .Z(n67469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54558_3_lut.init = 16'hcaca;
    LUT4 i54557_3_lut (.A(\hidden_outputs[0] [7]), .B(\hidden_outputs[1] [7]), 
         .C(n[0]), .Z(n67468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54557_3_lut.init = 16'hcaca;
    LUT4 i54555_3_lut (.A(\hidden_outputs[2] [6]), .B(\hidden_outputs[3] [6]), 
         .C(n[0]), .Z(n67466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54555_3_lut.init = 16'hcaca;
    LUT4 i54554_3_lut (.A(\hidden_outputs[0] [6]), .B(\hidden_outputs[1] [6]), 
         .C(n[0]), .Z(n67465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54554_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_57 (.A(\hidden_outputs[1] [0]), .B(n22568), .C(float_alu_c[0]), 
         .D(n70789), .Z(n23360)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_57.init = 16'hc088;
    LUT4 i2_4_lut_adj_58 (.A(n23360), .B(n10_adj_77), .C(\hidden_outputs[1] [0]), 
         .D(n2022[17]), .Z(n63188)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_58.init = 16'hfeee;
    LUT4 select_455_Select_21_i32_2_lut (.A(sram_output_B[21]), .B(n2022[31]), 
         .Z(n32_adj_106)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_21_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_59 (.A(\mlp_outputs[1] [21]), .B(n70809), .C(float_alu_c[21]), 
         .D(o[0]), .Z(n22802)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_59.init = 16'hc088;
    LUT4 i1_4_lut_adj_60 (.A(n32_adj_106), .B(n22802), .C(\mlp_outputs[1] [21]), 
         .D(n2022[39]), .Z(n66454)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_60.init = 16'hfeee;
    LUT4 select_455_Select_22_i32_2_lut (.A(sram_output_B[22]), .B(n2022[31]), 
         .Z(n32_adj_107)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_22_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_61 (.A(\mlp_outputs[1] [22]), .B(n70809), .C(float_alu_c[22]), 
         .D(o[0]), .Z(n23207)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_61.init = 16'hc088;
    LUT4 i1_4_lut_adj_62 (.A(n32_adj_107), .B(\mlp_outputs[1] [22]), .C(n23207), 
         .D(n2022[39]), .Z(n66298)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_62.init = 16'hfefa;
    PFUMX i54346 (.BLUT(n67255), .ALUT(n67256), .C0(h[1]), .Z(n67257));
    CCU2D add_4597_10 (.A0(\i[8] ), .B0(h[9]), .C0(GND_net), .D0(GND_net), 
          .A1(\i[9] ), .B1(h[10]), .C1(GND_net), .D1(GND_net), .CIN(n61480), 
          .COUT(n61481), .S0(n7729[8]), .S1(n7729[9]));
    defparam add_4597_10.INIT0 = 16'h5666;
    defparam add_4597_10.INIT1 = 16'h5666;
    defparam add_4597_10.INJECT1_0 = "NO";
    defparam add_4597_10.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(n2022[19]), .B(n2022[27]), .Z(n6_adj_108)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(n2022[23]), .B(n6_adj_108), .C(n2022[25]), .D(n2022[21]), 
         .Z(n66196)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    CCU2D add_4584_add_1_add_1_5 (.A0(n14054), .B0(numL[0]), .C0(n12), 
          .D0(n929), .A1(n14054), .B1(numL[0]), .C1(n12), .D1(n928), 
          .CIN(n61483), .COUT(n61484), .S0(n3[3]), .S1(n3[4]));
    defparam add_4584_add_1_add_1_5.INIT0 = 16'hfe00;
    defparam add_4584_add_1_add_1_5.INIT1 = 16'hfe00;
    defparam add_4584_add_1_add_1_5.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_5.INJECT1_1 = "NO";
    FD1S3AX No_Name_i1 (.D(\buf_x[83] ), .CK(clock), .Q(\buf_r[83] ));
    defparam No_Name_i1.GSR = "DISABLED";
    PFUMX i54349 (.BLUT(n67258), .ALUT(n67259), .C0(i[1]), .Z(n67260));
    LUT4 i2_2_lut_adj_63 (.A(n2082), .B(n66196), .Z(n6_adj_109)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_adj_63.init = 16'heeee;
    FD1P3AX temp_outputs_0__i0_i6 (.D(\hidden_outputs[0] [6]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [6]));
    defparam temp_outputs_0__i0_i6.GSR = "DISABLED";
    LUT4 i29161_4_lut (.A(n70822), .B(n2022[17]), .C(n6_adj_109), .D(n70846), 
         .Z(n40754)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i29161_4_lut.init = 16'haaa8;
    LUT4 select_450_Select_0_i10_2_lut (.A(sram_output_B[0]), .B(n2022[9]), 
         .Z(n10_adj_77)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_0_i10_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_64 (.A(n2022[49]), .B(n27496), .Z(n3756)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_64.init = 16'h2222;
    LUT4 i1_4_lut_adj_65 (.A(n73818), .B(n2082), .C(n27496), .D(n2022[49]), 
         .Z(n77)) /* synthesis lut_function=(!((B (C (D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_65.init = 16'h0a88;
    CCU2D equal_97_24 (.A0(i_c[31]), .B0(i_c[30]), .C0(i_c[29]), .D0(i_c[28]), 
          .A1(i_c[28]), .B1(i_c[27]), .C1(i_c[26]), .D1(i_c[25]), .CIN(n60973), 
          .COUT(n60974));
    defparam equal_97_24.INIT0 = 16'h8001;
    defparam equal_97_24.INIT1 = 16'h8001;
    defparam equal_97_24.INJECT1_0 = "YES";
    defparam equal_97_24.INJECT1_1 = "YES";
    LUT4 i1_2_lut_adj_66 (.A(n66196), .B(n2022[16]), .Z(n22568)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_66.init = 16'heeee;
    LUT4 i1_4_lut_adj_67 (.A(\hidden_outputs[0] [0]), .B(n22568), .C(float_alu_c[0]), 
         .D(n70791), .Z(n22748)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_67.init = 16'h88c0;
    FD1P3AX output_outputs_0__i0_i31 (.D(n66434), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [31]));
    defparam output_outputs_0__i0_i31.GSR = "DISABLED";
    CCU2D equal_97_0 (.A0(i_c[31]), .B0(n3921), .C0(GND_net), .D0(GND_net), 
          .A1(i[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n60973));
    defparam equal_97_0.INIT0 = 16'h9000;
    defparam equal_97_0.INIT1 = 16'haaaa;
    defparam equal_97_0.INJECT1_0 = "NO";
    defparam equal_97_0.INJECT1_1 = "YES";
    PFUMX i54355 (.BLUT(n67264), .ALUT(n67265), .C0(i[1]), .Z(n67266));
    LUT4 i2_4_lut_adj_68 (.A(n10_adj_77), .B(n22748), .C(\hidden_outputs[0] [0]), 
         .D(n2022[17]), .Z(n62956)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_68.init = 16'hfeee;
    CCU2D add_4584_add_1_add_1_11 (.A0(n14054), .B0(numL[0]), .C0(n12), 
          .D0(n923), .A1(n14054), .B1(numL[0]), .C1(n12), .D1(n922), 
          .CIN(n61486), .COUT(n61487), .S0(n3[9]), .S1(n3[10]));
    defparam add_4584_add_1_add_1_11.INIT0 = 16'hfe00;
    defparam add_4584_add_1_add_1_11.INIT1 = 16'hfe00;
    defparam add_4584_add_1_add_1_11.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_11.INJECT1_1 = "NO";
    LUT4 i2_3_lut (.A(mlp_ready), .B(\state[0] ), .C(mlp_mode), .Z(n63309)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut.init = 16'h0808;
    PFUMX i54358 (.BLUT(n67267), .ALUT(n67268), .C0(i[1]), .Z(n67269));
    LUT4 i54552_3_lut (.A(\hidden_outputs[2] [5]), .B(\hidden_outputs[3] [5]), 
         .C(n[0]), .Z(n67463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54552_3_lut.init = 16'hcaca;
    LUT4 i54551_3_lut (.A(\hidden_outputs[0] [5]), .B(\hidden_outputs[1] [5]), 
         .C(n[0]), .Z(n67462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54551_3_lut.init = 16'hcaca;
    PFUMX i54361 (.BLUT(n67270), .ALUT(n67271), .C0(i[1]), .Z(n67272));
    PFUMX i54364 (.BLUT(n67273), .ALUT(n67274), .C0(i[1]), .Z(n67275));
    PFUMX i54367 (.BLUT(n67276), .ALUT(n67277), .C0(i[1]), .Z(n67278));
    LUT4 select_455_Select_23_i32_2_lut (.A(sram_output_B[23]), .B(n2022[31]), 
         .Z(n32_adj_110)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_23_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_69 (.A(\mlp_outputs[1] [23]), .B(n70809), .C(float_alu_c[23]), 
         .D(o[0]), .Z(n23504)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_69.init = 16'hc088;
    LUT4 i1_4_lut_adj_70 (.A(n32_adj_110), .B(\mlp_outputs[1] [23]), .C(n23504), 
         .D(n2022[39]), .Z(n66340)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_70.init = 16'hfefa;
    LUT4 i1_4_lut_adj_71 (.A(\mlp_outputs[1] [0]), .B(n70809), .C(float_alu_c[0]), 
         .D(o[0]), .Z(n23351)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_71.init = 16'hc088;
    LUT4 i2_4_lut_adj_72 (.A(n23351), .B(n32_adj_111), .C(\mlp_outputs[1] [0]), 
         .D(n2022[39]), .Z(n63184)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_72.init = 16'hfeee;
    PFUMX i54370 (.BLUT(n67279), .ALUT(n67280), .C0(i[1]), .Z(n67281));
    FD1P3AX output_outputs_0__i0_i30 (.D(n66364), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [30]));
    defparam output_outputs_0__i0_i30.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i29 (.D(n62986), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [29]));
    defparam output_outputs_0__i0_i29.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i28 (.D(n66366), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [28]));
    defparam output_outputs_0__i0_i28.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i27 (.D(n63215), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [27]));
    defparam output_outputs_0__i0_i27.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i26 (.D(n62983), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [26]));
    defparam output_outputs_0__i0_i26.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i25 (.D(n66436), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [25]));
    defparam output_outputs_0__i0_i25.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i24 (.D(n63217), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [24]));
    defparam output_outputs_0__i0_i24.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i23 (.D(n62981), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [23]));
    defparam output_outputs_0__i0_i23.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i22 (.D(n66362), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [22]));
    defparam output_outputs_0__i0_i22.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i21 (.D(n66438), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [21]));
    defparam output_outputs_0__i0_i21.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i20 (.D(n63219), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [20]));
    defparam output_outputs_0__i0_i20.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i19 (.D(n66440), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [19]));
    defparam output_outputs_0__i0_i19.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i18 (.D(n62978), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [18]));
    defparam output_outputs_0__i0_i18.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i17 (.D(n63221), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [17]));
    defparam output_outputs_0__i0_i17.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i16 (.D(n62976), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [16]));
    defparam output_outputs_0__i0_i16.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i15 (.D(n66320), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [15]));
    defparam output_outputs_0__i0_i15.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i14 (.D(n66442), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [14]));
    defparam output_outputs_0__i0_i14.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i13 (.D(n63227), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [13]));
    defparam output_outputs_0__i0_i13.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i12 (.D(n63232), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [12]));
    defparam output_outputs_0__i0_i12.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i11 (.D(n66396), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [11]));
    defparam output_outputs_0__i0_i11.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i10 (.D(n66342), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [10]));
    defparam output_outputs_0__i0_i10.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i9 (.D(n66446), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [9]));
    defparam output_outputs_0__i0_i9.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i8 (.D(n63235), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [8]));
    defparam output_outputs_0__i0_i8.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i7 (.D(n62972), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [7]));
    defparam output_outputs_0__i0_i7.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i6 (.D(n66350), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [6]));
    defparam output_outputs_0__i0_i6.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i5 (.D(n66368), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [5]));
    defparam output_outputs_0__i0_i5.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i4 (.D(n62990), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [4]));
    defparam output_outputs_0__i0_i4.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i3 (.D(n63206), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [3]));
    defparam output_outputs_0__i0_i3.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i2 (.D(n63203), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [2]));
    defparam output_outputs_0__i0_i2.GSR = "DISABLED";
    FD1P3AX output_outputs_0__i0_i1 (.D(n63213), .SP(n23646), .CK(clock), 
            .Q(\mlp_outputs[0] [1]));
    defparam output_outputs_0__i0_i1.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i11 (.D(n63155), .SP(n23627), .CK(clock), .Q(sram_address_B[11]));
    defparam sram_addr_i0_i11.GSR = "DISABLED";
    PFUMX i54373 (.BLUT(n67282), .ALUT(n67283), .C0(i[1]), .Z(n67284));
    PFUMX i54376 (.BLUT(n67285), .ALUT(n67286), .C0(i[1]), .Z(n67287));
    LUT4 i55131_2_lut (.A(\float_alu_mode[2] ), .B(n1155), .Z(n124)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i55131_2_lut.init = 16'h1111;
    LUT4 i54549_3_lut (.A(\hidden_outputs[2] [4]), .B(\hidden_outputs[3] [4]), 
         .C(n[0]), .Z(n67460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54549_3_lut.init = 16'hcaca;
    LUT4 i54548_3_lut (.A(\hidden_outputs[0] [4]), .B(\hidden_outputs[1] [4]), 
         .C(n[0]), .Z(n67459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54548_3_lut.init = 16'hcaca;
    LUT4 i54546_3_lut (.A(\hidden_outputs[2] [3]), .B(\hidden_outputs[3] [3]), 
         .C(n[0]), .Z(n67457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54546_3_lut.init = 16'hcaca;
    LUT4 i54545_3_lut (.A(\hidden_outputs[0] [3]), .B(\hidden_outputs[1] [3]), 
         .C(n[0]), .Z(n67456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54545_3_lut.init = 16'hcaca;
    LUT4 i54543_3_lut (.A(\hidden_outputs[2] [2]), .B(\hidden_outputs[3] [2]), 
         .C(n[0]), .Z(n67454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54543_3_lut.init = 16'hcaca;
    LUT4 i54542_3_lut (.A(\hidden_outputs[0] [2]), .B(\hidden_outputs[1] [2]), 
         .C(n[0]), .Z(n67453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54542_3_lut.init = 16'hcaca;
    LUT4 i54540_3_lut (.A(\hidden_outputs[2] [1]), .B(\hidden_outputs[3] [1]), 
         .C(n[0]), .Z(n67451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54540_3_lut.init = 16'hcaca;
    FD1P3AX sram_addr_i0_i10 (.D(n63119), .SP(n23627), .CK(clock), .Q(sram_address_B[10]));
    defparam sram_addr_i0_i10.GSR = "DISABLED";
    LUT4 i54539_3_lut (.A(\hidden_outputs[0] [1]), .B(\hidden_outputs[1] [1]), 
         .C(n[0]), .Z(n67450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54539_3_lut.init = 16'hcaca;
    LUT4 i54537_3_lut (.A(\hidden_outputs[2] [31]), .B(\hidden_outputs[3] [31]), 
         .C(h[0]), .Z(n67448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54537_3_lut.init = 16'hcaca;
    LUT4 i54536_3_lut (.A(\hidden_outputs[0] [31]), .B(\hidden_outputs[1] [31]), 
         .C(h[0]), .Z(n67447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54536_3_lut.init = 16'hcaca;
    LUT4 i54534_3_lut (.A(\hidden_outputs[2] [30]), .B(\hidden_outputs[3] [30]), 
         .C(h[0]), .Z(n67445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54534_3_lut.init = 16'hcaca;
    LUT4 i54533_3_lut (.A(\hidden_outputs[0] [30]), .B(\hidden_outputs[1] [30]), 
         .C(h[0]), .Z(n67444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54533_3_lut.init = 16'hcaca;
    PFUMX i54379 (.BLUT(n67288), .ALUT(n67289), .C0(i[1]), .Z(n67290));
    LUT4 i54531_3_lut (.A(\hidden_outputs[2] [29]), .B(\hidden_outputs[3] [29]), 
         .C(h[0]), .Z(n67442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54531_3_lut.init = 16'hcaca;
    LUT4 i54530_3_lut (.A(\hidden_outputs[0] [29]), .B(\hidden_outputs[1] [29]), 
         .C(h[0]), .Z(n67441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54530_3_lut.init = 16'hcaca;
    LUT4 i54528_3_lut (.A(\hidden_outputs[2] [28]), .B(\hidden_outputs[3] [28]), 
         .C(h[0]), .Z(n67439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54528_3_lut.init = 16'hcaca;
    LUT4 i54527_3_lut (.A(\hidden_outputs[0] [28]), .B(\hidden_outputs[1] [28]), 
         .C(h[0]), .Z(n67438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54527_3_lut.init = 16'hcaca;
    LUT4 i54525_3_lut (.A(\hidden_outputs[2] [27]), .B(\hidden_outputs[3] [27]), 
         .C(h[0]), .Z(n67436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54525_3_lut.init = 16'hcaca;
    LUT4 i54524_3_lut (.A(\hidden_outputs[0] [27]), .B(\hidden_outputs[1] [27]), 
         .C(h[0]), .Z(n67435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54524_3_lut.init = 16'hcaca;
    LUT4 i54522_3_lut (.A(\hidden_outputs[2] [26]), .B(\hidden_outputs[3] [26]), 
         .C(h[0]), .Z(n67433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54522_3_lut.init = 16'hcaca;
    LUT4 i54521_3_lut (.A(\hidden_outputs[0] [26]), .B(\hidden_outputs[1] [26]), 
         .C(h[0]), .Z(n67432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54521_3_lut.init = 16'hcaca;
    LUT4 i54519_3_lut (.A(\hidden_outputs[2] [25]), .B(\hidden_outputs[3] [25]), 
         .C(h[0]), .Z(n67430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54519_3_lut.init = 16'hcaca;
    LUT4 i54518_3_lut (.A(\hidden_outputs[0] [25]), .B(\hidden_outputs[1] [25]), 
         .C(h[0]), .Z(n67429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54518_3_lut.init = 16'hcaca;
    LUT4 i54516_3_lut (.A(\hidden_outputs[2] [24]), .B(\hidden_outputs[3] [24]), 
         .C(h[0]), .Z(n67427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54516_3_lut.init = 16'hcaca;
    LUT4 i54515_3_lut (.A(\hidden_outputs[0] [24]), .B(\hidden_outputs[1] [24]), 
         .C(h[0]), .Z(n67426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54515_3_lut.init = 16'hcaca;
    FD1P3DX float_alu_mode_i0_i2 (.D(n23975), .SP(n27939), .CK(clock), 
            .CD(SDA_c), .Q(\float_alu_mode[2] ));
    defparam float_alu_mode_i0_i2.GSR = "DISABLED";
    LUT4 i1_3_lut (.A(n2022[12]), .B(n70822), .C(n2022[34]), .Z(n4593)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut.init = 16'hc8c8;
    FD1P3IX addr_4653__i31 (.D(n134_adj_408[31]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[31]));
    defparam addr_4653__i31.GSR = "DISABLED";
    FD1P3IX addr_4653__i27 (.D(n134_adj_408[27]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[27]));
    defparam addr_4653__i27.GSR = "DISABLED";
    FD1P3IX addr_4653__i28 (.D(n134_adj_408[28]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[28]));
    defparam addr_4653__i28.GSR = "DISABLED";
    FD1P3IX addr_4653__i29 (.D(n134_adj_408[29]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[29]));
    defparam addr_4653__i29.GSR = "DISABLED";
    FD1P3IX addr_4653__i26 (.D(n134_adj_408[26]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[26]));
    defparam addr_4653__i26.GSR = "DISABLED";
    FD1P3IX addr_4653__i30 (.D(n134_adj_408[30]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[30]));
    defparam addr_4653__i30.GSR = "DISABLED";
    FD1P3IX addr_4653__i22 (.D(n134_adj_408[22]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[22]));
    defparam addr_4653__i22.GSR = "DISABLED";
    FD1P3IX addr_4653__i16 (.D(n134_adj_408[16]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[16]));
    defparam addr_4653__i16.GSR = "DISABLED";
    FD1P3IX addr_4653__i23 (.D(n134_adj_408[23]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[23]));
    defparam addr_4653__i23.GSR = "DISABLED";
    FD1P3IX addr_4653__i17 (.D(n134_adj_408[17]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[17]));
    defparam addr_4653__i17.GSR = "DISABLED";
    FD1P3IX addr_4653__i12 (.D(n134_adj_408[12]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[12]));
    defparam addr_4653__i12.GSR = "DISABLED";
    FD1P3IX addr_4653__i18 (.D(n134_adj_408[18]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[18]));
    defparam addr_4653__i18.GSR = "DISABLED";
    FD1P3IX addr_4653__i24 (.D(n134_adj_408[24]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[24]));
    defparam addr_4653__i24.GSR = "DISABLED";
    FD1P3IX addr_4653__i19 (.D(n134_adj_408[19]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[19]));
    defparam addr_4653__i19.GSR = "DISABLED";
    FD1P3IX addr_4653__i13 (.D(n134_adj_408[13]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[13]));
    defparam addr_4653__i13.GSR = "DISABLED";
    FD1P3IX addr_4653__i20 (.D(n134_adj_408[20]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[20]));
    defparam addr_4653__i20.GSR = "DISABLED";
    FD1P3IX addr_4653__i14 (.D(n134_adj_408[14]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[14]));
    defparam addr_4653__i14.GSR = "DISABLED";
    FD1P3IX addr_4653__i15 (.D(n134_adj_408[15]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[15]));
    defparam addr_4653__i15.GSR = "DISABLED";
    FD1P3IX addr_4653__i21 (.D(n134_adj_408[21]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[21]));
    defparam addr_4653__i21.GSR = "DISABLED";
    FD1P3IX addr_4653__i25 (.D(n134_adj_408[25]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[25]));
    defparam addr_4653__i25.GSR = "DISABLED";
    FD1P3IX addr_4653__i3 (.D(n134_adj_408[3]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[3]));
    defparam addr_4653__i3.GSR = "DISABLED";
    FD1P3IX addr_4653__i9 (.D(n134_adj_408[9]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[9]));
    defparam addr_4653__i9.GSR = "DISABLED";
    FD1P3IX addr_4653__i4 (.D(n134_adj_408[4]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[4]));
    defparam addr_4653__i4.GSR = "DISABLED";
    FD1P3IX numL_4656__i30 (.D(n134_adj_407[30]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[30]));
    defparam numL_4656__i30.GSR = "DISABLED";
    FD1P3IX addr_4653__i5 (.D(n134_adj_408[5]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[5]));
    defparam addr_4653__i5.GSR = "DISABLED";
    FD1P3IX addr_4653__i10 (.D(n134_adj_408[10]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[10]));
    defparam addr_4653__i10.GSR = "DISABLED";
    FD1P3IX addr_4653__i6 (.D(n134_adj_408[6]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[6]));
    defparam addr_4653__i6.GSR = "DISABLED";
    FD1P3IX numL_4656__i31 (.D(n134_adj_407[31]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[31]));
    defparam numL_4656__i31.GSR = "DISABLED";
    FD1P3IX addr_4653__i7 (.D(n134_adj_408[7]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[7]));
    defparam addr_4653__i7.GSR = "DISABLED";
    FD1P3IX addr_4653__i1 (.D(n134_adj_408[1]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[1]));
    defparam addr_4653__i1.GSR = "DISABLED";
    FD1P3IX addr_4653__i2 (.D(n134_adj_408[2]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[2]));
    defparam addr_4653__i2.GSR = "DISABLED";
    FD1P3IX addr_4653__i8 (.D(n134_adj_408[8]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[8]));
    defparam addr_4653__i8.GSR = "DISABLED";
    FD1P3IX addr_4653__i11 (.D(n134_adj_408[11]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[11]));
    defparam addr_4653__i11.GSR = "DISABLED";
    FD1P3IX numL_4656__i28 (.D(n134_adj_407[28]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[28]));
    defparam numL_4656__i28.GSR = "DISABLED";
    FD1P3IX numL_4656__i29 (.D(n134_adj_407[29]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[29]));
    defparam numL_4656__i29.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i9 (.D(n63158), .SP(n23627), .CK(clock), .Q(sram_address_B[9]));
    defparam sram_addr_i0_i9.GSR = "DISABLED";
    FD1P3IX numL_4656__i17 (.D(n134_adj_407[17]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[17]));
    defparam numL_4656__i17.GSR = "DISABLED";
    FD1P3IX numL_4656__i24 (.D(n134_adj_407[24]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[24]));
    defparam numL_4656__i24.GSR = "DISABLED";
    FD1P3IX numL_4656__i10 (.D(n134_adj_407[10]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[10]));
    defparam numL_4656__i10.GSR = "DISABLED";
    FD1P3IX numL_4656__i18 (.D(n134_adj_407[18]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[18]));
    defparam numL_4656__i18.GSR = "DISABLED";
    FD1P3IX numL_4656__i25 (.D(n134_adj_407[25]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[25]));
    defparam numL_4656__i25.GSR = "DISABLED";
    FD1P3IX numL_4656__i11 (.D(n134_adj_407[11]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[11]));
    defparam numL_4656__i11.GSR = "DISABLED";
    FD1P3IX numL_4656__i19 (.D(n134_adj_407[19]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[19]));
    defparam numL_4656__i19.GSR = "DISABLED";
    FD1P3IX numL_4656__i5 (.D(n134_adj_407[5]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[5]));
    defparam numL_4656__i5.GSR = "DISABLED";
    FD1P3IX numL_4656__i12 (.D(n134_adj_407[12]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[12]));
    defparam numL_4656__i12.GSR = "DISABLED";
    FD1P3IX numL_4656__i20 (.D(n134_adj_407[20]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[20]));
    defparam numL_4656__i20.GSR = "DISABLED";
    FD1P3IX numL_4656__i26 (.D(n134_adj_407[26]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[26]));
    defparam numL_4656__i26.GSR = "DISABLED";
    FD1P3IX numL_4656__i13 (.D(n134_adj_407[13]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[13]));
    defparam numL_4656__i13.GSR = "DISABLED";
    FD1P3IX numL_4656__i21 (.D(n134_adj_407[21]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[21]));
    defparam numL_4656__i21.GSR = "DISABLED";
    FD1P3IX numL_4656__i6 (.D(n134_adj_407[6]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[6]));
    defparam numL_4656__i6.GSR = "DISABLED";
    FD1P3IX numL_4656__i14 (.D(n134_adj_407[14]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[14]));
    defparam numL_4656__i14.GSR = "DISABLED";
    FD1P3IX numL_4656__i22 (.D(n134_adj_407[22]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[22]));
    defparam numL_4656__i22.GSR = "DISABLED";
    FD1P3IX numL_4656__i7 (.D(n134_adj_407[7]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[7]));
    defparam numL_4656__i7.GSR = "DISABLED";
    FD1P3IX numL_4656__i15 (.D(n134_adj_407[15]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[15]));
    defparam numL_4656__i15.GSR = "DISABLED";
    FD1P3IX numL_4656__i8 (.D(n134_adj_407[8]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[8]));
    defparam numL_4656__i8.GSR = "DISABLED";
    FD1P3IX numL_4656__i9 (.D(n134_adj_407[9]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[9]));
    defparam numL_4656__i9.GSR = "DISABLED";
    FD1P3IX numL_4656__i16 (.D(n134_adj_407[16]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[16]));
    defparam numL_4656__i16.GSR = "DISABLED";
    FD1P3IX numL_4656__i23 (.D(n134_adj_407[23]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[23]));
    defparam numL_4656__i23.GSR = "DISABLED";
    FD1P3IX numL_4656__i27 (.D(n134_adj_407[27]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[27]));
    defparam numL_4656__i27.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i8 (.D(n63163), .SP(n23627), .CK(clock), .Q(sram_address_B[8]));
    defparam sram_addr_i0_i8.GSR = "DISABLED";
    FD1P3IX h_4657__i30 (.D(n134[30]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[30]));
    defparam h_4657__i30.GSR = "DISABLED";
    FD1P3IX h_4657__i15 (.D(n134[15]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[15]));
    defparam h_4657__i15.GSR = "DISABLED";
    FD1P3IX h_4657__i31 (.D(n134[31]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[31]));
    defparam h_4657__i31.GSR = "DISABLED";
    FD1P3IX h_4657__i16 (.D(n134[16]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[16]));
    defparam h_4657__i16.GSR = "DISABLED";
    FD1P3IX h_4657__i17 (.D(n134[17]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[17]));
    defparam h_4657__i17.GSR = "DISABLED";
    FD1P3IX numL_4656__i1 (.D(n134_adj_407[1]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(n14054));
    defparam numL_4656__i1.GSR = "DISABLED";
    FD1P3IX h_4657__i18 (.D(n134[18]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[18]));
    defparam h_4657__i18.GSR = "DISABLED";
    FD1P3IX h_4657__i19 (.D(n134[19]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[19]));
    defparam h_4657__i19.GSR = "DISABLED";
    FD1P3IX h_4657__i20 (.D(n134[20]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[20]));
    defparam h_4657__i20.GSR = "DISABLED";
    FD1P3IX numL_4656__i2 (.D(n134_adj_407[2]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[2]));
    defparam numL_4656__i2.GSR = "DISABLED";
    FD1P3IX h_4657__i21 (.D(n134[21]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[21]));
    defparam h_4657__i21.GSR = "DISABLED";
    FD1P3IX n_4659__i30 (.D(n134_adj_403[30]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[30]));
    defparam n_4659__i30.GSR = "DISABLED";
    FD1P3IX h_4657__i22 (.D(n134[22]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[22]));
    defparam h_4657__i22.GSR = "DISABLED";
    FD1P3IX n_4659__i31 (.D(n134_adj_403[31]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[31]));
    defparam n_4659__i31.GSR = "DISABLED";
    FD1P3IX h_4657__i1 (.D(n134[1]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[1]));
    defparam h_4657__i1.GSR = "DISABLED";
    FD1P3IX h_4657__i23 (.D(n134[23]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[23]));
    defparam h_4657__i23.GSR = "DISABLED";
    FD1P3IX h_4657__i2 (.D(n134[2]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[2]));
    defparam h_4657__i2.GSR = "DISABLED";
    FD1P3IX h_4657__i3 (.D(n134[3]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[3]));
    defparam h_4657__i3.GSR = "DISABLED";
    FD1P3IX h_4657__i4 (.D(n134[4]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[4]));
    defparam h_4657__i4.GSR = "DISABLED";
    FD1P3IX h_4657__i24 (.D(n134[24]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[24]));
    defparam h_4657__i24.GSR = "DISABLED";
    FD1P3IX numL_4656__i3 (.D(n134_adj_407[3]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[3]));
    defparam numL_4656__i3.GSR = "DISABLED";
    FD1P3IX h_4657__i25 (.D(n134[25]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[25]));
    defparam h_4657__i25.GSR = "DISABLED";
    FD1P3IX h_4657__i5 (.D(n134[5]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[5]));
    defparam h_4657__i5.GSR = "DISABLED";
    FD1P3IX h_4657__i26 (.D(n134[26]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[26]));
    defparam h_4657__i26.GSR = "DISABLED";
    FD1P3IX h_4657__i6 (.D(n134[6]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[6]));
    defparam h_4657__i6.GSR = "DISABLED";
    FD1P3IX h_4657__i7 (.D(n134[7]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[7]));
    defparam h_4657__i7.GSR = "DISABLED";
    FD1P3IX h_4657__i27 (.D(n134[27]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[27]));
    defparam h_4657__i27.GSR = "DISABLED";
    FD1P3IX h_4657__i8 (.D(n134[8]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[8]));
    defparam h_4657__i8.GSR = "DISABLED";
    FD1P3IX h_4657__i9 (.D(n134[9]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[9]));
    defparam h_4657__i9.GSR = "DISABLED";
    FD1P3IX h_4657__i10 (.D(n134[10]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[10]));
    defparam h_4657__i10.GSR = "DISABLED";
    FD1P3IX h_4657__i28 (.D(n134[28]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[28]));
    defparam h_4657__i28.GSR = "DISABLED";
    FD1P3IX h_4657__i11 (.D(n134[11]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[11]));
    defparam h_4657__i11.GSR = "DISABLED";
    FD1P3IX h_4657__i12 (.D(n134[12]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[12]));
    defparam h_4657__i12.GSR = "DISABLED";
    FD1P3IX h_4657__i13 (.D(n134[13]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[13]));
    defparam h_4657__i13.GSR = "DISABLED";
    FD1P3IX h_4657__i14 (.D(n134[14]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[14]));
    defparam h_4657__i14.GSR = "DISABLED";
    FD1P3IX h_4657__i29 (.D(n134[29]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[29]));
    defparam h_4657__i29.GSR = "DISABLED";
    FD1P3IX numL_4656__i4 (.D(n134_adj_407[4]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[4]));
    defparam numL_4656__i4.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i7 (.D(n63164), .SP(n23627), .CK(clock), .Q(sram_address_B[7]));
    defparam sram_addr_i0_i7.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i6 (.D(n63167), .SP(n23627), .CK(clock), .Q(sram_address_B[6]));
    defparam sram_addr_i0_i6.GSR = "DISABLED";
    FD1P3DX state_FSM__i49 (.D(n66556), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2036));
    defparam state_FSM__i49.GSR = "DISABLED";
    FD1P3DX state_FSM__i48 (.D(n2022[48]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[49]));
    defparam state_FSM__i48.GSR = "DISABLED";
    FD1P3DX state_FSM__i47 (.D(n2022[47]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[48]));
    defparam state_FSM__i47.GSR = "DISABLED";
    FD1P3DX state_FSM__i46 (.D(n2022[46]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[47]));
    defparam state_FSM__i46.GSR = "DISABLED";
    FD1P3DX state_FSM__i45 (.D(n2022[45]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[46]));
    defparam state_FSM__i45.GSR = "DISABLED";
    FD1P3DX state_FSM__i44 (.D(n2022[44]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[45]));
    defparam state_FSM__i44.GSR = "DISABLED";
    FD1P3DX state_FSM__i43 (.D(n2022[43]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[44]));
    defparam state_FSM__i43.GSR = "DISABLED";
    FD1P3DX state_FSM__i42 (.D(n2022[42]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[43]));
    defparam state_FSM__i42.GSR = "DISABLED";
    FD1P3DX state_FSM__i41 (.D(n2022[41]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[42]));
    defparam state_FSM__i41.GSR = "DISABLED";
    FD1P3DX state_FSM__i40 (.D(n2022[40]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[41]));
    defparam state_FSM__i40.GSR = "DISABLED";
    FD1P3DX state_FSM__i39 (.D(n2022[39]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[40]));
    defparam state_FSM__i39.GSR = "DISABLED";
    FD1P3DX state_FSM__i38 (.D(n2284), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[39]));
    defparam state_FSM__i38.GSR = "DISABLED";
    FD1P3DX state_FSM__i37 (.D(n2022[37]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[38]));
    defparam state_FSM__i37.GSR = "DISABLED";
    FD1P3DX state_FSM__i36 (.D(n2050), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[37]));
    defparam state_FSM__i36.GSR = "DISABLED";
    FD1P3DX state_FSM__i35 (.D(n2022[35]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2050));
    defparam state_FSM__i35.GSR = "DISABLED";
    FD1P3DX state_FSM__i34 (.D(n2022[34]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[35]));
    defparam state_FSM__i34.GSR = "DISABLED";
    FD1P3DX state_FSM__i33 (.D(n2022[33]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[34]));
    defparam state_FSM__i33.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i5 (.D(n63255), .SP(n23627), .CK(clock), .Q(sram_address_B[5]));
    defparam sram_addr_i0_i5.GSR = "DISABLED";
    FD1P3DX state_FSM__i32 (.D(n2022[32]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[33]));
    defparam state_FSM__i32.GSR = "DISABLED";
    FD1P3DX state_FSM__i31 (.D(n2277), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[32]));
    defparam state_FSM__i31.GSR = "DISABLED";
    FD1P3DX state_FSM__i30 (.D(n2022[30]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[31]));
    defparam state_FSM__i30.GSR = "DISABLED";
    FD1P3DX state_FSM__i29 (.D(n2022[29]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[30]));
    defparam state_FSM__i29.GSR = "DISABLED";
    FD1P3DX state_FSM__i28 (.D(n2272), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[29]));
    defparam state_FSM__i28.GSR = "DISABLED";
    FD1P3DX state_FSM__i27 (.D(n2269), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[28]));
    defparam state_FSM__i27.GSR = "DISABLED";
    FD1P3DX state_FSM__i26 (.D(n2022[26]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[27]));
    defparam state_FSM__i26.GSR = "DISABLED";
    FD1P3DX state_FSM__i25 (.D(n2022[25]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[26]));
    defparam state_FSM__i25.GSR = "DISABLED";
    FD1P3DX state_FSM__i24 (.D(n2022[24]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[25]));
    defparam state_FSM__i24.GSR = "DISABLED";
    FD1P3DX state_FSM__i23 (.D(n2022[23]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[24]));
    defparam state_FSM__i23.GSR = "DISABLED";
    FD1P3DX state_FSM__i22 (.D(n2022[22]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[23]));
    defparam state_FSM__i22.GSR = "DISABLED";
    FD1P3DX state_FSM__i21 (.D(n2022[21]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[22]));
    defparam state_FSM__i21.GSR = "DISABLED";
    FD1P3DX state_FSM__i20 (.D(n2022[20]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[21]));
    defparam state_FSM__i20.GSR = "DISABLED";
    FD1P3DX state_FSM__i19 (.D(n2022[19]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[20]));
    defparam state_FSM__i19.GSR = "DISABLED";
    FD1P3DX state_FSM__i18 (.D(n2022[18]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[19]));
    defparam state_FSM__i18.GSR = "DISABLED";
    FD1P3DX state_FSM__i17 (.D(n2022[17]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[18]));
    defparam state_FSM__i17.GSR = "DISABLED";
    FD1P3DX state_FSM__i16 (.D(n70701), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[17]));
    defparam state_FSM__i16.GSR = "DISABLED";
    FD1P3DX state_FSM__i15 (.D(n2022[15]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[16]));
    defparam state_FSM__i15.GSR = "DISABLED";
    FD1P3DX state_FSM__i14 (.D(n2072), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[15]));
    defparam state_FSM__i14.GSR = "DISABLED";
    FD1P3DX state_FSM__i13 (.D(n2022[13]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2072));
    defparam state_FSM__i13.GSR = "DISABLED";
    FD1P3DX state_FSM__i12 (.D(n2022[12]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[13]));
    defparam state_FSM__i12.GSR = "DISABLED";
    FD1P3DX state_FSM__i11 (.D(n2022[11]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[12]));
    defparam state_FSM__i11.GSR = "DISABLED";
    FD1P3DX state_FSM__i10 (.D(n2022[10]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[11]));
    defparam state_FSM__i10.GSR = "DISABLED";
    FD1P3DX state_FSM__i9 (.D(n2251), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[10]));
    defparam state_FSM__i9.GSR = "DISABLED";
    FD1P3DX state_FSM__i8 (.D(n2022[8]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[9]));
    defparam state_FSM__i8.GSR = "DISABLED";
    FD1P3DX state_FSM__i7 (.D(n2022[7]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[8]));
    defparam state_FSM__i7.GSR = "DISABLED";
    FD1P3DX state_FSM__i6 (.D(n63041), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[7]));
    defparam state_FSM__i6.GSR = "DISABLED";
    FD1P3DX state_FSM__i5 (.D(n2242), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2082));
    defparam state_FSM__i5.GSR = "DISABLED";
    FD1P3DX state_FSM__i4 (.D(n2084), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[3]));
    defparam state_FSM__i4.GSR = "DISABLED";
    FD1P3DX state_FSM__i3 (.D(n2022[1]), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2084));
    defparam state_FSM__i3.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i4 (.D(n63238), .SP(n23627), .CK(clock), .Q(sram_address_B[4]));
    defparam sram_addr_i0_i4.GSR = "DISABLED";
    FD1P3DX state_FSM__i2 (.D(n2239), .SP(n70816), .CK(clock), .CD(SDA_c), 
            .Q(n2022[1]));
    defparam state_FSM__i2.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i3 (.D(n63138), .SP(n23627), .CK(clock), .Q(sram_address_B[3]));
    defparam sram_addr_i0_i3.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i2 (.D(n63135), .SP(n23627), .CK(clock), .Q(sram_address_B[2]));
    defparam sram_addr_i0_i2.GSR = "DISABLED";
    FD1P3AX sram_addr_i0_i1 (.D(n63018), .SP(n23627), .CK(clock), .Q(sram_address_B[1]));
    defparam sram_addr_i0_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n22276), .B(n70768), .C(n70822), .D(n70858), 
         .Z(n23664)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0e0;
    PFUMX i54382 (.BLUT(n67291), .ALUT(n67292), .C0(i[1]), .Z(n67293));
    PFUMX i54385 (.BLUT(n67294), .ALUT(n67295), .C0(i[1]), .Z(n67296));
    FD1P3AX f_i0_i31 (.D(float_alu_c[31]), .SP(n4617), .CK(clock), .Q(f[31]));
    defparam f_i0_i31.GSR = "DISABLED";
    FD1P3AX f_i0_i30 (.D(float_alu_c[30]), .SP(n4617), .CK(clock), .Q(f[30]));
    defparam f_i0_i30.GSR = "DISABLED";
    FD1P3AX f_i0_i29 (.D(float_alu_c[29]), .SP(n4617), .CK(clock), .Q(f[29]));
    defparam f_i0_i29.GSR = "DISABLED";
    FD1P3AX f_i0_i28 (.D(float_alu_c[28]), .SP(n4617), .CK(clock), .Q(f[28]));
    defparam f_i0_i28.GSR = "DISABLED";
    FD1P3AX f_i0_i27 (.D(float_alu_c[27]), .SP(n4617), .CK(clock), .Q(f[27]));
    defparam f_i0_i27.GSR = "DISABLED";
    FD1P3AX f_i0_i26 (.D(float_alu_c[26]), .SP(n4617), .CK(clock), .Q(f[26]));
    defparam f_i0_i26.GSR = "DISABLED";
    FD1P3AX f_i0_i25 (.D(float_alu_c[25]), .SP(n4617), .CK(clock), .Q(f[25]));
    defparam f_i0_i25.GSR = "DISABLED";
    FD1P3AX f_i0_i24 (.D(float_alu_c[24]), .SP(n4617), .CK(clock), .Q(f[24]));
    defparam f_i0_i24.GSR = "DISABLED";
    FD1P3AX f_i0_i23 (.D(float_alu_c[23]), .SP(n4617), .CK(clock), .Q(f[23]));
    defparam f_i0_i23.GSR = "DISABLED";
    FD1P3AX f_i0_i22 (.D(float_alu_c[22]), .SP(n4617), .CK(clock), .Q(f[22]));
    defparam f_i0_i22.GSR = "DISABLED";
    FD1P3AX f_i0_i21 (.D(float_alu_c[21]), .SP(n4617), .CK(clock), .Q(f[21]));
    defparam f_i0_i21.GSR = "DISABLED";
    FD1P3AX f_i0_i20 (.D(float_alu_c[20]), .SP(n4617), .CK(clock), .Q(f[20]));
    defparam f_i0_i20.GSR = "DISABLED";
    FD1P3AX f_i0_i19 (.D(float_alu_c[19]), .SP(n4617), .CK(clock), .Q(f[19]));
    defparam f_i0_i19.GSR = "DISABLED";
    FD1P3AX f_i0_i18 (.D(float_alu_c[18]), .SP(n4617), .CK(clock), .Q(f[18]));
    defparam f_i0_i18.GSR = "DISABLED";
    FD1P3AX f_i0_i17 (.D(float_alu_c[17]), .SP(n4617), .CK(clock), .Q(f[17]));
    defparam f_i0_i17.GSR = "DISABLED";
    FD1P3AX f_i0_i16 (.D(float_alu_c[16]), .SP(n4617), .CK(clock), .Q(f[16]));
    defparam f_i0_i16.GSR = "DISABLED";
    FD1P3AX f_i0_i15 (.D(float_alu_c[15]), .SP(n4617), .CK(clock), .Q(f[15]));
    defparam f_i0_i15.GSR = "DISABLED";
    FD1P3AX f_i0_i14 (.D(float_alu_c[14]), .SP(n4617), .CK(clock), .Q(f[14]));
    defparam f_i0_i14.GSR = "DISABLED";
    FD1P3AX f_i0_i13 (.D(float_alu_c[13]), .SP(n4617), .CK(clock), .Q(f[13]));
    defparam f_i0_i13.GSR = "DISABLED";
    FD1P3AX f_i0_i12 (.D(float_alu_c[12]), .SP(n4617), .CK(clock), .Q(f[12]));
    defparam f_i0_i12.GSR = "DISABLED";
    FD1P3AX f_i0_i11 (.D(float_alu_c[11]), .SP(n4617), .CK(clock), .Q(f[11]));
    defparam f_i0_i11.GSR = "DISABLED";
    FD1P3AX f_i0_i10 (.D(float_alu_c[10]), .SP(n4617), .CK(clock), .Q(f[10]));
    defparam f_i0_i10.GSR = "DISABLED";
    FD1P3AX f_i0_i9 (.D(float_alu_c[9]), .SP(n4617), .CK(clock), .Q(f[9]));
    defparam f_i0_i9.GSR = "DISABLED";
    FD1P3AX f_i0_i8 (.D(float_alu_c[8]), .SP(n4617), .CK(clock), .Q(f[8]));
    defparam f_i0_i8.GSR = "DISABLED";
    FD1P3AX f_i0_i7 (.D(float_alu_c[7]), .SP(n4617), .CK(clock), .Q(f[7]));
    defparam f_i0_i7.GSR = "DISABLED";
    FD1P3AX f_i0_i6 (.D(float_alu_c[6]), .SP(n4617), .CK(clock), .Q(f[6]));
    defparam f_i0_i6.GSR = "DISABLED";
    FD1P3AX f_i0_i5 (.D(float_alu_c[5]), .SP(n4617), .CK(clock), .Q(f[5]));
    defparam f_i0_i5.GSR = "DISABLED";
    FD1P3AX f_i0_i4 (.D(float_alu_c[4]), .SP(n4617), .CK(clock), .Q(f[4]));
    defparam f_i0_i4.GSR = "DISABLED";
    FD1P3AX f_i0_i3 (.D(float_alu_c[3]), .SP(n4617), .CK(clock), .Q(f[3]));
    defparam f_i0_i3.GSR = "DISABLED";
    FD1P3AX f_i0_i2 (.D(float_alu_c[2]), .SP(n4617), .CK(clock), .Q(f[2]));
    defparam f_i0_i2.GSR = "DISABLED";
    FD1P3AX f_i0_i1 (.D(float_alu_c[1]), .SP(n4617), .CK(clock), .Q(f[1]));
    defparam f_i0_i1.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i31 (.D(\hidden_outputs[0] [31]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [31]));
    defparam temp_outputs_0__i0_i31.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i30 (.D(\hidden_outputs[0] [30]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [30]));
    defparam temp_outputs_0__i0_i30.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i29 (.D(\hidden_outputs[0] [29]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [29]));
    defparam temp_outputs_0__i0_i29.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i28 (.D(\hidden_outputs[0] [28]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [28]));
    defparam temp_outputs_0__i0_i28.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i27 (.D(\hidden_outputs[0] [27]), .SP(n73808), 
            .CK(clock), .Q(\temp_outputs[0] [27]));
    defparam temp_outputs_0__i0_i27.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i26 (.D(\hidden_outputs[0] [26]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [26]));
    defparam temp_outputs_0__i0_i26.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i25 (.D(\hidden_outputs[0] [25]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [25]));
    defparam temp_outputs_0__i0_i25.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i24 (.D(\hidden_outputs[0] [24]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [24]));
    defparam temp_outputs_0__i0_i24.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i23 (.D(\hidden_outputs[0] [23]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [23]));
    defparam temp_outputs_0__i0_i23.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i22 (.D(\hidden_outputs[0] [22]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [22]));
    defparam temp_outputs_0__i0_i22.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i21 (.D(\hidden_outputs[0] [21]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [21]));
    defparam temp_outputs_0__i0_i21.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i20 (.D(\hidden_outputs[0] [20]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [20]));
    defparam temp_outputs_0__i0_i20.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i19 (.D(\hidden_outputs[0] [19]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [19]));
    defparam temp_outputs_0__i0_i19.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i18 (.D(\hidden_outputs[0] [18]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [18]));
    defparam temp_outputs_0__i0_i18.GSR = "DISABLED";
    FD1P3AX temp_outputs_0__i0_i17 (.D(\hidden_outputs[0] [17]), .SP(n4923), 
            .CK(clock), .Q(\temp_outputs[0] [17]));
    defparam temp_outputs_0__i0_i17.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i1 (.D(n62897), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [1]));
    defparam hidden_outputs_0__i0_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_743_3_lut_4_lut (.A(n70786), .B(n66671), .C(numL[31]), 
         .D(n14054), .Z(n70713)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i1_2_lut_rep_743_3_lut_4_lut.init = 16'hf0f1;
    PFUMX i54388 (.BLUT(n67297), .ALUT(n67298), .C0(i[1]), .Z(n67299));
    PFUMX i54391 (.BLUT(n67300), .ALUT(n67301), .C0(i[1]), .Z(n67302));
    PFUMX i54394 (.BLUT(n67303), .ALUT(n67304), .C0(i[1]), .Z(n67305));
    PFUMX i54397 (.BLUT(n67306), .ALUT(n67307), .C0(i[1]), .Z(n67308));
    LUT4 i2_2_lut_rep_753_3_lut (.A(n70786), .B(n66671), .C(n14054), .Z(n70723)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_2_lut_rep_753_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(n70786), .B(n66671), .C(numL[31]), .Z(n12)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    PFUMX i54400 (.BLUT(n67309), .ALUT(n67310), .C0(i[1]), .Z(n67311));
    PFUMX i54403 (.BLUT(n67312), .ALUT(n67313), .C0(i[1]), .Z(n67314));
    PFUMX i54406 (.BLUT(n67315), .ALUT(n67316), .C0(i[1]), .Z(n67317));
    PFUMX i54409 (.BLUT(n67318), .ALUT(n67319), .C0(i[1]), .Z(n67320));
    PFUMX i54412 (.BLUT(n67321), .ALUT(n67322), .C0(i[1]), .Z(n67323));
    PFUMX i54415 (.BLUT(n67324), .ALUT(n67325), .C0(i[1]), .Z(n67326));
    LUT4 n70822_bdd_3_lut (.A(n70822), .B(n2022[9]), .C(n2022[16]), .Z(n23968)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam n70822_bdd_3_lut.init = 16'h0808;
    PFUMX i54418 (.BLUT(n67327), .ALUT(n67328), .C0(i[1]), .Z(n67329));
    PFUMX i54421 (.BLUT(n67330), .ALUT(n67331), .C0(i[1]), .Z(n67332));
    PFUMX i54424 (.BLUT(n67333), .ALUT(n67334), .C0(i[1]), .Z(n67335));
    PFUMX i54427 (.BLUT(n67336), .ALUT(n67337), .C0(i[1]), .Z(n67338));
    PFUMX i54430 (.BLUT(n67339), .ALUT(n67340), .C0(i[1]), .Z(n67341));
    PFUMX i54433 (.BLUT(n67342), .ALUT(n67343), .C0(i[1]), .Z(n67344));
    PFUMX i54436 (.BLUT(n67345), .ALUT(n67346), .C0(i[1]), .Z(n67347));
    PFUMX i54439 (.BLUT(n67348), .ALUT(n67349), .C0(i[1]), .Z(n67350));
    FD1P3JX float_alu_b_i0_i28 (.D(n63159), .SP(n23664), .PD(n63295), 
            .CK(clock), .Q(float_alu_b[28]));
    defparam float_alu_b_i0_i28.GSR = "DISABLED";
    FD1P3JX float_alu_b_i0_i24 (.D(n63254), .SP(n23664), .PD(n63295), 
            .CK(clock), .Q(float_alu_b[24]));
    defparam float_alu_b_i0_i24.GSR = "DISABLED";
    FD1P3IX i_4655__i31 (.D(n134_adj_409[31]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[31]));
    defparam i_4655__i31.GSR = "DISABLED";
    FD1P3IX i_4655__i30 (.D(n134_adj_409[30]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[30]));
    defparam i_4655__i30.GSR = "DISABLED";
    FD1P3IX i_4655__i29 (.D(n134_adj_409[29]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[29]));
    defparam i_4655__i29.GSR = "DISABLED";
    FD1P3IX i_4655__i28 (.D(n134_adj_409[28]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[28]));
    defparam i_4655__i28.GSR = "DISABLED";
    PFUMX i54442 (.BLUT(n67351), .ALUT(n67352), .C0(i[1]), .Z(n67353));
    PFUMX i54445 (.BLUT(n67354), .ALUT(n67355), .C0(i[1]), .Z(n67356));
    PFUMX i54448 (.BLUT(n67357), .ALUT(n67358), .C0(h[1]), .Z(n67359));
    PFUMX i54451 (.BLUT(n67360), .ALUT(n67361), .C0(h[1]), .Z(n67362));
    FD1P3IX i_4655__i27 (.D(n134_adj_409[27]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[27]));
    defparam i_4655__i27.GSR = "DISABLED";
    FD1P3IX i_4655__i26 (.D(n134_adj_409[26]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[26]));
    defparam i_4655__i26.GSR = "DISABLED";
    LUT4 i54513_3_lut (.A(\hidden_outputs[2] [23]), .B(\hidden_outputs[3] [23]), 
         .C(h[0]), .Z(n67424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54513_3_lut.init = 16'hcaca;
    LUT4 i54512_3_lut (.A(\hidden_outputs[0] [23]), .B(\hidden_outputs[1] [23]), 
         .C(h[0]), .Z(n67423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54512_3_lut.init = 16'hcaca;
    LUT4 i54510_3_lut (.A(\hidden_outputs[2] [22]), .B(\hidden_outputs[3] [22]), 
         .C(h[0]), .Z(n67421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54510_3_lut.init = 16'hcaca;
    LUT4 i54509_3_lut (.A(\hidden_outputs[0] [22]), .B(\hidden_outputs[1] [22]), 
         .C(h[0]), .Z(n67420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54509_3_lut.init = 16'hcaca;
    LUT4 i54507_3_lut (.A(\hidden_outputs[2] [21]), .B(\hidden_outputs[3] [21]), 
         .C(h[0]), .Z(n67418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54507_3_lut.init = 16'hcaca;
    LUT4 i54506_3_lut (.A(\hidden_outputs[0] [21]), .B(\hidden_outputs[1] [21]), 
         .C(h[0]), .Z(n67417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54506_3_lut.init = 16'hcaca;
    LUT4 i54504_3_lut (.A(\hidden_outputs[2] [20]), .B(\hidden_outputs[3] [20]), 
         .C(h[0]), .Z(n67415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54504_3_lut.init = 16'hcaca;
    LUT4 i54503_3_lut (.A(\hidden_outputs[0] [20]), .B(\hidden_outputs[1] [20]), 
         .C(h[0]), .Z(n67414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54503_3_lut.init = 16'hcaca;
    FD1P3IX i_4655__i25 (.D(n134_adj_409[25]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[25]));
    defparam i_4655__i25.GSR = "DISABLED";
    LUT4 i54501_3_lut (.A(\hidden_outputs[2] [19]), .B(\hidden_outputs[3] [19]), 
         .C(h[0]), .Z(n67412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54501_3_lut.init = 16'hcaca;
    LUT4 i54500_3_lut (.A(\hidden_outputs[0] [19]), .B(\hidden_outputs[1] [19]), 
         .C(h[0]), .Z(n67411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54500_3_lut.init = 16'hcaca;
    LUT4 i54498_3_lut (.A(\hidden_outputs[2] [18]), .B(\hidden_outputs[3] [18]), 
         .C(h[0]), .Z(n67409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54498_3_lut.init = 16'hcaca;
    LUT4 i54497_3_lut (.A(\hidden_outputs[0] [18]), .B(\hidden_outputs[1] [18]), 
         .C(h[0]), .Z(n67408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54497_3_lut.init = 16'hcaca;
    LUT4 i54495_3_lut (.A(\hidden_outputs[2] [17]), .B(\hidden_outputs[3] [17]), 
         .C(h[0]), .Z(n67406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54495_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_rep_908 (.A(n70731), .B(n14054), .C(n4613), 
         .D(numL[31]), .Z(n73806)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_rep_908.init = 16'hf010;
    LUT4 i12567_2_lut_3_lut_3_lut (.A(n2269), .B(n70822), .C(n27496), 
         .D(n2022[49]), .Z(n24257)) /* synthesis lut_function=(!(((D)+!B)+!A)) */ ;
    defparam i12567_2_lut_3_lut_3_lut.init = 16'h0088;
    LUT4 i54494_3_lut (.A(\hidden_outputs[0] [17]), .B(\hidden_outputs[1] [17]), 
         .C(h[0]), .Z(n67405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54494_3_lut.init = 16'hcaca;
    PFUMX i54454 (.BLUT(n67363), .ALUT(n67364), .C0(h[1]), .Z(n67365));
    PFUMX i54457 (.BLUT(n67366), .ALUT(n67367), .C0(h[1]), .Z(n67368));
    PFUMX i54460 (.BLUT(n67369), .ALUT(n67370), .C0(h[1]), .Z(n67371));
    LUT4 i54492_3_lut (.A(\hidden_outputs[2] [16]), .B(\hidden_outputs[3] [16]), 
         .C(h[0]), .Z(n67403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54492_3_lut.init = 16'hcaca;
    LUT4 i54491_3_lut (.A(\hidden_outputs[0] [16]), .B(\hidden_outputs[1] [16]), 
         .C(h[0]), .Z(n67402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54491_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_73 (.A(\hidden_outputs[4] [31]), .B(n22568), .C(float_alu_c[31]), 
         .D(n70783), .Z(n22733)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_73.init = 16'hc088;
    LUT4 i2_4_lut_adj_74 (.A(n10_adj_182), .B(n22733), .C(n1582), .D(n2022[17]), 
         .Z(n62951)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_74.init = 16'hfeee;
    LUT4 i1_4_lut_adj_75 (.A(\hidden_outputs[4] [30]), .B(n22568), .C(float_alu_c[30]), 
         .D(n70783), .Z(n23282)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_75.init = 16'hc088;
    PFUMX i54463 (.BLUT(n67372), .ALUT(n67373), .C0(h[1]), .Z(n67374));
    PFUMX i54466 (.BLUT(n67375), .ALUT(n67376), .C0(h[1]), .Z(n67377));
    PFUMX i54469 (.BLUT(n67378), .ALUT(n67379), .C0(h[1]), .Z(n67380));
    LUT4 i2_4_lut_adj_76 (.A(n23282), .B(n10_adj_183), .C(\hidden_outputs[4] [30]), 
         .D(n2022[17]), .Z(n63065)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_76.init = 16'hfeee;
    LUT4 i1_4_lut_adj_77 (.A(\hidden_outputs[4] [29]), .B(n22568), .C(float_alu_c[29]), 
         .D(n70783), .Z(n23369)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_77.init = 16'hc088;
    FD1P3IX i_4655__i24 (.D(n134_adj_409[24]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[24]));
    defparam i_4655__i24.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_78 (.A(n10_adj_185), .B(\hidden_outputs[4] [29]), 
         .C(n23369), .D(n2022[17]), .Z(n66384)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_78.init = 16'hfefa;
    LUT4 i1_4_lut_adj_79 (.A(\hidden_outputs[4] [28]), .B(n22568), .C(float_alu_c[28]), 
         .D(n70783), .Z(n22739)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_79.init = 16'hc088;
    LUT4 i2_4_lut_adj_80 (.A(n10_adj_186), .B(n22739), .C(\hidden_outputs[4] [28]), 
         .D(n2022[17]), .Z(n62953)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_80.init = 16'hfeee;
    LUT4 i1_4_lut_adj_81 (.A(\hidden_outputs[4] [27]), .B(n22568), .C(float_alu_c[27]), 
         .D(n70783), .Z(n22913)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_81.init = 16'hc088;
    LUT4 i1_4_lut_adj_82 (.A(n10_adj_187), .B(n22913), .C(\hidden_outputs[4] [27]), 
         .D(n2022[17]), .Z(n66408)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_82.init = 16'hfeee;
    LUT4 i1_4_lut_adj_83 (.A(\hidden_outputs[4] [26]), .B(n22568), .C(float_alu_c[26]), 
         .D(n70783), .Z(n22545)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_83.init = 16'hc088;
    LUT4 i1_4_lut_adj_84 (.A(n10_adj_188), .B(\hidden_outputs[4] [26]), 
         .C(n22545), .D(n2022[17]), .Z(n66326)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_84.init = 16'hfefa;
    LUT4 i1_4_lut_adj_85 (.A(\hidden_outputs[4] [25]), .B(n22568), .C(float_alu_c[25]), 
         .D(n70783), .Z(n23261)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_85.init = 16'hc088;
    LUT4 i1_4_lut_adj_86 (.A(n10_adj_189), .B(\hidden_outputs[4] [25]), 
         .C(n23261), .D(n2022[17]), .Z(n66498)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_86.init = 16'hfefa;
    LUT4 i1_4_lut_adj_87 (.A(\hidden_outputs[4] [24]), .B(n22568), .C(float_alu_c[24]), 
         .D(n70783), .Z(n23447)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_87.init = 16'hc088;
    LUT4 i1_4_lut_adj_88 (.A(n10_adj_190), .B(\hidden_outputs[4] [24]), 
         .C(n23447), .D(n2022[17]), .Z(n66360)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_88.init = 16'hfefa;
    PFUMX i54472 (.BLUT(n67381), .ALUT(n67382), .C0(h[1]), .Z(n67383));
    LUT4 i1_4_lut_adj_89 (.A(\hidden_outputs[4] [23]), .B(n22568), .C(float_alu_c[23]), 
         .D(n70783), .Z(n23366)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_89.init = 16'hc088;
    LUT4 i2_4_lut_adj_90 (.A(n23366), .B(n10_adj_191), .C(\hidden_outputs[4] [23]), 
         .D(n2022[17]), .Z(n63190)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_90.init = 16'hfeee;
    LUT4 i1_4_lut_adj_91 (.A(\hidden_outputs[4] [22]), .B(n22568), .C(float_alu_c[22]), 
         .D(n70783), .Z(n22916)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_91.init = 16'hc088;
    LUT4 i2_4_lut_adj_92 (.A(n10_adj_192), .B(n22916), .C(\hidden_outputs[4] [22]), 
         .D(n2022[17]), .Z(n63014)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_92.init = 16'hfeee;
    LUT4 i1_4_lut_adj_93 (.A(\hidden_outputs[4] [21]), .B(n22568), .C(float_alu_c[21]), 
         .D(n70783), .Z(n22928)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_93.init = 16'hc088;
    LUT4 i1_4_lut_adj_94 (.A(n10_adj_193), .B(n22928), .C(\hidden_outputs[4] [21]), 
         .D(n2022[17]), .Z(n66318)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_94.init = 16'hfeee;
    LUT4 i1_4_lut_adj_95 (.A(\hidden_outputs[4] [20]), .B(n22568), .C(float_alu_c[20]), 
         .D(n70783), .Z(n23192)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_95.init = 16'hc088;
    PFUMX i54475 (.BLUT(n67384), .ALUT(n67385), .C0(h[1]), .Z(n67386));
    PFUMX i54478 (.BLUT(n67387), .ALUT(n67388), .C0(h[1]), .Z(n67389));
    LUT4 i1_4_lut_adj_96 (.A(n10_adj_194), .B(\hidden_outputs[4] [20]), 
         .C(n23192), .D(n2022[17]), .Z(n66302)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_96.init = 16'hfefa;
    LUT4 i1_4_lut_adj_97 (.A(\hidden_outputs[4] [19]), .B(n22568), .C(float_alu_c[19]), 
         .D(n70783), .Z(n22943)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_97.init = 16'hc088;
    LUT4 i1_4_lut_adj_98 (.A(n10_adj_195), .B(n22943), .C(\hidden_outputs[4] [19]), 
         .D(n2022[17]), .Z(n66270)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_98.init = 16'hfeee;
    LUT4 i1_4_lut_adj_99 (.A(\hidden_outputs[4] [18]), .B(n22568), .C(float_alu_c[18]), 
         .D(n70783), .Z(n23354)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_99.init = 16'hc088;
    LUT4 i1_4_lut_adj_100 (.A(n10_adj_196), .B(\hidden_outputs[4] [18]), 
         .C(n23354), .D(n2022[17]), .Z(n66388)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_100.init = 16'hfefa;
    LUT4 i1_4_lut_adj_101 (.A(\hidden_outputs[4] [17]), .B(n22568), .C(float_alu_c[17]), 
         .D(n70783), .Z(n23519)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_101.init = 16'hc088;
    FD1P3IX i_4655__i23 (.D(n134_adj_409[23]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[23]));
    defparam i_4655__i23.GSR = "DISABLED";
    FD1P3IX i_4655__i22 (.D(n134_adj_409[22]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[22]));
    defparam i_4655__i22.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_102 (.A(n10_adj_199), .B(\hidden_outputs[4] [17]), 
         .C(n23519), .D(n2022[17]), .Z(n66330)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_102.init = 16'hfefa;
    FD1P3IX i_4655__i21 (.D(n134_adj_409[21]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[21]));
    defparam i_4655__i21.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_103 (.A(\hidden_outputs[4] [16]), .B(n22568), .C(float_alu_c[16]), 
         .D(n70783), .Z(n22946)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_103.init = 16'hc088;
    FD1P3IX i_4655__i20 (.D(n134_adj_409[20]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[20]));
    defparam i_4655__i20.GSR = "DISABLED";
    FD1P3IX i_4655__i19 (.D(n134_adj_409[19]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[19]));
    defparam i_4655__i19.GSR = "DISABLED";
    FD1P3IX i_4655__i18 (.D(n134_adj_409[18]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[18]));
    defparam i_4655__i18.GSR = "DISABLED";
    FD1P3IX i_4655__i17 (.D(n134_adj_409[17]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[17]));
    defparam i_4655__i17.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_104 (.A(n10_adj_205), .B(n22946), .C(\hidden_outputs[4] [16]), 
         .D(n2022[17]), .Z(n66398)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_104.init = 16'hfeee;
    LUT4 i1_4_lut_adj_105 (.A(\hidden_outputs[4] [15]), .B(n22568), .C(float_alu_c[15]), 
         .D(n70783), .Z(n22940)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_105.init = 16'hc088;
    FD1P3IX i_4655__i16 (.D(n134_adj_409[16]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[16]));
    defparam i_4655__i16.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_106 (.A(n10_adj_207), .B(n22940), .C(\hidden_outputs[4] [15]), 
         .D(n2022[17]), .Z(n66276)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_106.init = 16'hfeee;
    LUT4 i1_4_lut_adj_107 (.A(\hidden_outputs[4] [14]), .B(n22568), .C(float_alu_c[14]), 
         .D(n70783), .Z(n22563)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_107.init = 16'hc088;
    FD1P3IX i_4655__i15 (.D(n134_adj_409[15]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[15]));
    defparam i_4655__i15.GSR = "DISABLED";
    FD1P3IX i_4655__i14 (.D(n134_adj_409[14]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[14]));
    defparam i_4655__i14.GSR = "DISABLED";
    FD1P3IX i_4655__i13 (.D(n134_adj_409[13]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i_c[13]));
    defparam i_4655__i13.GSR = "DISABLED";
    FD1P3IX i_4655__i12 (.D(n134_adj_409[12]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[12] ));
    defparam i_4655__i12.GSR = "DISABLED";
    FD1P3IX i_4655__i11 (.D(n134_adj_409[11]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[11] ));
    defparam i_4655__i11.GSR = "DISABLED";
    FD1P3IX i_4655__i10 (.D(n134_adj_409[10]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i[10]));
    defparam i_4655__i10.GSR = "DISABLED";
    FD1P3IX i_4655__i9 (.D(n134_adj_409[9]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[9] ));
    defparam i_4655__i9.GSR = "DISABLED";
    FD1P3IX i_4655__i8 (.D(n134_adj_409[8]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[8] ));
    defparam i_4655__i8.GSR = "DISABLED";
    FD1P3IX i_4655__i7 (.D(n134_adj_409[7]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[7] ));
    defparam i_4655__i7.GSR = "DISABLED";
    FD1P3IX i_4655__i6 (.D(n134_adj_409[6]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[6] ));
    defparam i_4655__i6.GSR = "DISABLED";
    FD1P3IX i_4655__i5 (.D(n134_adj_409[5]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[5] ));
    defparam i_4655__i5.GSR = "DISABLED";
    FD1P3IX i_4655__i4 (.D(n134_adj_409[4]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[4] ));
    defparam i_4655__i4.GSR = "DISABLED";
    FD1P3IX i_4655__i3 (.D(n134_adj_409[3]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(\i[3] ));
    defparam i_4655__i3.GSR = "DISABLED";
    FD1P3IX i_4655__i2 (.D(n134_adj_409[2]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i[2]));
    defparam i_4655__i2.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_108 (.A(n10_adj_222), .B(n22563), .C(\hidden_outputs[4] [14]), 
         .D(n2022[17]), .Z(n66536)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_108.init = 16'hfeee;
    FD1P3IX i_4655__i1 (.D(n134_adj_409[1]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i[1]));
    defparam i_4655__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_109 (.A(\hidden_outputs[4] [13]), .B(n22568), .C(float_alu_c[13]), 
         .D(n70783), .Z(n22760)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_109.init = 16'hc088;
    LUT4 i1_4_lut_adj_110 (.A(n10_adj_224), .B(n22760), .C(\hidden_outputs[4] [13]), 
         .D(n2022[17]), .Z(n66462)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_110.init = 16'hfeee;
    LUT4 i1_4_lut_adj_111 (.A(\hidden_outputs[4] [12]), .B(n22568), .C(float_alu_c[12]), 
         .D(n70783), .Z(n22551)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_111.init = 16'hc088;
    LUT4 i1_4_lut_adj_112 (.A(n10_adj_225), .B(\hidden_outputs[4] [12]), 
         .C(n22551), .D(n2022[17]), .Z(n66268)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_112.init = 16'hfefa;
    LUT4 i1_4_lut_adj_113 (.A(\hidden_outputs[4] [11]), .B(n22568), .C(float_alu_c[11]), 
         .D(n70783), .Z(n22778)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_113.init = 16'hc088;
    LUT4 i1_4_lut_adj_114 (.A(n10_adj_226), .B(\hidden_outputs[4] [11]), 
         .C(n22778), .D(n2022[17]), .Z(n66450)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_114.init = 16'hfefa;
    LUT4 i1_4_lut_adj_115 (.A(\hidden_outputs[4] [10]), .B(n22568), .C(float_alu_c[10]), 
         .D(n70783), .Z(n23198)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_115.init = 16'hc088;
    LUT4 i1_4_lut_adj_116 (.A(n10_adj_227), .B(\hidden_outputs[4] [10]), 
         .C(n23198), .D(n2022[17]), .Z(n66286)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_116.init = 16'hfefa;
    LUT4 i1_4_lut_adj_117 (.A(\hidden_outputs[4] [9]), .B(n22568), .C(float_alu_c[9]), 
         .D(n70783), .Z(n23138)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_117.init = 16'hc088;
    LUT4 i1_4_lut_adj_118 (.A(n10_adj_228), .B(\hidden_outputs[4] [9]), 
         .C(n23138), .D(n2022[17]), .Z(n66424)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_118.init = 16'hfefa;
    LUT4 i1_4_lut_adj_119 (.A(\hidden_outputs[4] [8]), .B(n22568), .C(float_alu_c[8]), 
         .D(n70783), .Z(n22811)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_119.init = 16'hc088;
    LUT4 i1_4_lut_adj_120 (.A(n10_adj_229), .B(\hidden_outputs[4] [8]), 
         .C(n22811), .D(n2022[17]), .Z(n66550)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_120.init = 16'hfefa;
    LUT4 i1_4_lut_adj_121 (.A(\hidden_outputs[4] [7]), .B(n22568), .C(float_alu_c[7]), 
         .D(n70783), .Z(n23531)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_121.init = 16'hc088;
    LUT4 i1_4_lut_adj_122 (.A(n10_adj_230), .B(\hidden_outputs[4] [7]), 
         .C(n23531), .D(n2022[17]), .Z(n66328)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_122.init = 16'hfefa;
    LUT4 i1_4_lut_adj_123 (.A(\hidden_outputs[4] [6]), .B(n22568), .C(float_alu_c[6]), 
         .D(n70783), .Z(n23318)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_123.init = 16'hc088;
    LUT4 i1_4_lut_adj_124 (.A(n10_adj_231), .B(\hidden_outputs[4] [6]), 
         .C(n23318), .D(n2022[17]), .Z(n66546)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_124.init = 16'hfefa;
    LUT4 i1_4_lut_adj_125 (.A(\hidden_outputs[4] [5]), .B(n22568), .C(float_alu_c[5]), 
         .D(n70783), .Z(n22577)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_125.init = 16'hc088;
    LUT4 i2_4_lut_adj_126 (.A(n10_adj_232), .B(n22577), .C(\hidden_outputs[4] [5]), 
         .D(n2022[17]), .Z(n62864)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_126.init = 16'hfeee;
    LUT4 i1_4_lut_adj_127 (.A(\hidden_outputs[4] [4]), .B(n22568), .C(float_alu_c[4]), 
         .D(n70783), .Z(n22625)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_127.init = 16'hc088;
    LUT4 i1_4_lut_adj_128 (.A(n10_adj_233), .B(n22625), .C(\hidden_outputs[4] [4]), 
         .D(n2022[17]), .Z(n66516)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_128.init = 16'hfeee;
    LUT4 i1_4_lut_adj_129 (.A(\hidden_outputs[4] [3]), .B(n22568), .C(float_alu_c[3]), 
         .D(n70783), .Z(n23492)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_129.init = 16'hc088;
    LUT4 i1_4_lut_adj_130 (.A(n10_adj_234), .B(\hidden_outputs[4] [3]), 
         .C(n23492), .D(n2022[17]), .Z(n66344)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_130.init = 16'hfefa;
    LUT4 i1_4_lut_adj_131 (.A(\hidden_outputs[4] [2]), .B(n22568), .C(float_alu_c[2]), 
         .D(n70783), .Z(n22736)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_131.init = 16'hc088;
    LUT4 i1_4_lut_adj_132 (.A(n10_adj_235), .B(n22736), .C(\hidden_outputs[4] [2]), 
         .D(n2022[17]), .Z(n66470)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_132.init = 16'hfeee;
    LUT4 i1_4_lut_adj_133 (.A(\hidden_outputs[4] [1]), .B(n22568), .C(float_alu_c[1]), 
         .D(n70783), .Z(n23273)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_133.init = 16'hc088;
    LUT4 i1_4_lut_adj_134 (.A(n10_adj_236), .B(\hidden_outputs[4] [1]), 
         .C(n23273), .D(n2022[17]), .Z(n66282)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_134.init = 16'hfefa;
    LUT4 i1_4_lut_rep_904 (.A(n2269), .B(n70822), .C(n27496), .D(n2022[49]), 
         .Z(n73800)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_rep_904.init = 16'hc088;
    LUT4 mux_75_Mux_31_i7_4_lut (.A(n67269), .B(\temp_outputs[4] [31]), 
         .C(i[2]), .D(n17802), .Z(n1028[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_31_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i32_3_lut (.A(n1028[31]), .B(n1027[31]), .C(n70712), .Z(n1061[31])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i32_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_135 (.A(f[31]), .B(n2448[31]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_237)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_135.init = 16'heca0;
    LUT4 select_460_Select_31_i16_2_lut (.A(e[31]), .B(n2022[15]), .Z(n16_adj_238)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_31_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_136 (.A(n17745), .B(n8_adj_237), .C(n1061[31]), 
         .D(n2022[13]), .Z(n10_adj_239)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_136.init = 16'hfeee;
    LUT4 mux_220_Mux_31_i7_4_lut (.A(n67542), .B(\hidden_outputs[4] [31]), 
         .C(n[2]), .D(n70842), .Z(n3742[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_31_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_137 (.A(n3742[31]), .B(n10_adj_239), .C(n16_adj_238), 
         .D(n2022[35]), .Z(n63021)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_137.init = 16'hfefc;
    LUT4 mux_75_Mux_30_i7_4_lut (.A(n67272), .B(\temp_outputs[4] [30]), 
         .C(i[2]), .D(n17802), .Z(n1028[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_30_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i31_3_lut (.A(n1028[30]), .B(n1027[30]), .C(n70712), .Z(n1061[30])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i31_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_138 (.A(f[30]), .B(n2448[30]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_240)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_138.init = 16'heca0;
    LUT4 select_460_Select_30_i16_2_lut (.A(e[30]), .B(n2022[15]), .Z(n16_adj_241)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_30_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_139 (.A(n17726), .B(n8_adj_240), .C(n1061[30]), 
         .D(n2022[13]), .Z(n10_adj_242)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_139.init = 16'hfeee;
    LUT4 mux_220_Mux_30_i7_4_lut (.A(n67539), .B(\hidden_outputs[4] [30]), 
         .C(n[2]), .D(n70842), .Z(n3742[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_30_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_140 (.A(n3742[30]), .B(n10_adj_242), .C(n16_adj_241), 
         .D(n2022[35]), .Z(n63151)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_140.init = 16'hfefc;
    LUT4 mux_75_Mux_29_i7_4_lut (.A(n67275), .B(\temp_outputs[4] [29]), 
         .C(i[2]), .D(n17802), .Z(n1028[29])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_29_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i30_3_lut (.A(n1028[29]), .B(n1027[29]), .C(n70712), .Z(n1061[29])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i30_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_141 (.A(n1061[29]), .B(n4478[29]), .C(n2022[13]), 
         .D(n70843), .Z(n8_adj_243)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_141.init = 16'heca0;
    LUT4 select_460_Select_29_i36_4_lut (.A(n67536), .B(n2022[35]), .C(n6_adj_244), 
         .D(n[2]), .Z(n36_adj_245)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam select_460_Select_29_i36_4_lut.init = 16'hc088;
    LUT4 i4_4_lut_adj_142 (.A(n22931), .B(n8_adj_243), .C(e[29]), .D(n2022[15]), 
         .Z(n10_adj_246)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_142.init = 16'hfeee;
    LUT4 select_460_Select_29_i38_2_lut (.A(f[29]), .B(n2022[37]), .Z(n38_adj_247)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_29_i38_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_143 (.A(n22424), .B(n38_adj_247), .C(n10_adj_246), 
         .D(n36_adj_245), .Z(n66484)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_143.init = 16'hfffe;
    LUT4 mux_75_Mux_27_i7_4_lut (.A(n67281), .B(\temp_outputs[4] [27]), 
         .C(i[2]), .D(n17802), .Z(n1028[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_27_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i28_3_lut (.A(n1028[27]), .B(n1027[27]), .C(n70712), .Z(n1061[27])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i28_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_144 (.A(n1061[27]), .B(n4478[27]), .C(n2022[13]), 
         .D(n70843), .Z(n8_adj_248)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_144.init = 16'heca0;
    LUT4 select_460_Select_27_i36_4_lut (.A(n67530), .B(n2022[35]), .C(n6_adj_249), 
         .D(n[2]), .Z(n36_adj_250)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam select_460_Select_27_i36_4_lut.init = 16'hc088;
    LUT4 i4_4_lut_adj_145 (.A(n22934), .B(n8_adj_248), .C(e[27]), .D(n2022[15]), 
         .Z(n10_adj_251)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_145.init = 16'hfeee;
    LUT4 select_460_Select_27_i38_2_lut (.A(f[27]), .B(n2022[37]), .Z(n38_adj_252)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_27_i38_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_146 (.A(n22424), .B(n38_adj_252), .C(n10_adj_251), 
         .D(n36_adj_250), .Z(n66310)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_146.init = 16'hfffe;
    PFUMX i54481 (.BLUT(n67390), .ALUT(n67391), .C0(h[1]), .Z(n67392));
    LUT4 mux_141_Mux_26_i7_4_lut (.A(n67434), .B(\hidden_outputs[4] [26]), 
         .C(h[2]), .D(n70861), .Z(n2448[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_26_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_26_i1_3_lut (.A(\mlp_outputs[0] [26]), .B(\mlp_outputs[1] [26]), 
         .C(o[0]), .Z(n4478[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_26_i1_3_lut.init = 16'hcaca;
    LUT4 mux_75_Mux_26_i7_4_lut (.A(n67284), .B(\temp_outputs[4] [26]), 
         .C(i[2]), .D(n17802), .Z(n1028[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_26_i7_4_lut.init = 16'h0aca;
    LUT4 i1_3_lut_rep_746_4_lut (.A(n70858), .B(n70736), .C(n70859), .D(n70822), 
         .Z(n70716)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_rep_746_4_lut.init = 16'hfe00;
    LUT4 mux_76_i27_3_lut (.A(n1028[26]), .B(n1027[26]), .C(n70712), .Z(n1061[26])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i27_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_147 (.A(n1061[26]), .B(n4478[26]), .C(n2022[13]), 
         .D(n70843), .Z(n8_adj_253)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_147.init = 16'heca0;
    LUT4 select_460_Select_26_i36_4_lut (.A(n67527), .B(n2022[35]), .C(n6_adj_254), 
         .D(n[2]), .Z(n36_adj_255)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam select_460_Select_26_i36_4_lut.init = 16'hc088;
    LUT4 i4_4_lut_adj_148 (.A(n22925), .B(n8_adj_253), .C(e[26]), .D(n2022[15]), 
         .Z(n10_adj_256)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_148.init = 16'hfeee;
    LUT4 select_460_Select_26_i38_2_lut (.A(f[26]), .B(n2022[37]), .Z(n38_adj_257)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_26_i38_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_149 (.A(n22424), .B(n38_adj_257), .C(n10_adj_256), 
         .D(n36_adj_255), .Z(n66412)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_149.init = 16'hfffe;
    LUT4 i1_2_lut_rep_754 (.A(n2022[49]), .B(n27496), .Z(n70724)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_754.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_150 (.A(n70731), .B(n14054), .C(n2022[28]), 
         .D(numL[31]), .Z(n35)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_150.init = 16'hf010;
    LUT4 mux_75_Mux_25_i7_4_lut (.A(n67287), .B(\temp_outputs[4] [25]), 
         .C(i[2]), .D(n17802), .Z(n1028[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_25_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i26_3_lut (.A(n1028[25]), .B(n1027[25]), .C(n70712), .Z(n1061[25])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i26_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_4_lut_adj_151 (.A(n70731), .B(n14054), .C(n4613), 
         .D(numL[31]), .Z(n4923)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_151.init = 16'hf010;
    LUT4 i2_4_lut_adj_152 (.A(n1061[25]), .B(n4478[25]), .C(n2022[13]), 
         .D(n70843), .Z(n8_adj_258)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_152.init = 16'heca0;
    LUT4 select_460_Select_25_i36_4_lut (.A(n67524), .B(n2022[35]), .C(n6_adj_259), 
         .D(n[2]), .Z(n36_adj_260)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam select_460_Select_25_i36_4_lut.init = 16'hc088;
    LUT4 i4_4_lut_adj_153 (.A(n22922), .B(n8_adj_258), .C(e[25]), .D(n2022[15]), 
         .Z(n10_adj_261)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_153.init = 16'hfeee;
    LUT4 select_460_Select_25_i38_2_lut (.A(f[25]), .B(n2022[37]), .Z(n38_adj_262)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_25_i38_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_154 (.A(n22424), .B(n38_adj_262), .C(n10_adj_261), 
         .D(n36_adj_260), .Z(n66404)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_154.init = 16'hfffe;
    LUT4 select_455_Select_24_i32_2_lut (.A(sram_output_B[24]), .B(n2022[31]), 
         .Z(n32_adj_263)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_24_i32_2_lut.init = 16'h8888;
    PFUMX i54484 (.BLUT(n67393), .ALUT(n67394), .C0(h[1]), .Z(n67395));
    LUT4 mux_220_Mux_23_i7_4_lut (.A(n67518), .B(\hidden_outputs[4] [23]), 
         .C(n[2]), .D(n70842), .Z(n3742[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_23_i7_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_155 (.A(\mlp_outputs[1] [24]), .B(n70809), .C(float_alu_c[24]), 
         .D(o[0]), .Z(n22805)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_155.init = 16'hc088;
    LUT4 i3_3_lut_rep_742_4_lut (.A(n70731), .B(n14054), .C(numL[31]), 
         .D(numL[0]), .Z(n70712)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_742_4_lut.init = 16'hfffe;
    LUT4 mux_75_Mux_23_i7_4_lut (.A(n67293), .B(\temp_outputs[4] [23]), 
         .C(i[2]), .D(n17802), .Z(n1028[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_23_i7_4_lut.init = 16'h0aca;
    LUT4 i2_4_lut_adj_156 (.A(n32_adj_263), .B(n22805), .C(\mlp_outputs[1] [24]), 
         .D(n2022[39]), .Z(n62969)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_156.init = 16'hfeee;
    LUT4 i3_4_lut_adj_157 (.A(f[23]), .B(n3742[23]), .C(n2022[37]), .D(n2022[35]), 
         .Z(n10_adj_264)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_157.init = 16'heca0;
    LUT4 mux_76_i24_3_lut (.A(n1028[23]), .B(n1027[23]), .C(n70712), .Z(n1061[23])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i24_3_lut.init = 16'hacac;
    LUT4 select_460_Select_23_i16_2_lut (.A(e[23]), .B(n2022[15]), .Z(n16_adj_265)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_23_i16_2_lut.init = 16'h8888;
    LUT4 i5_4_lut_adj_158 (.A(n1061[23]), .B(n10_adj_264), .C(n17644), 
         .D(n2022[13]), .Z(n12_adj_266)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_158.init = 16'hfefc;
    LUT4 i6_4_lut (.A(n22424), .B(n12_adj_266), .C(n22919), .D(n16_adj_265), 
         .Z(n63015)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 mux_75_Mux_22_i7_4_lut (.A(n67296), .B(\temp_outputs[4] [22]), 
         .C(i[2]), .D(n17802), .Z(n1028[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_22_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i23_3_lut (.A(n1028[22]), .B(n1027[22]), .C(n70712), .Z(n1061[22])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i23_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_159 (.A(f[22]), .B(n2448[22]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_267)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_159.init = 16'heca0;
    LUT4 select_460_Select_22_i16_2_lut (.A(e[22]), .B(n2022[15]), .Z(n16_adj_268)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_22_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_160 (.A(n17638), .B(n8_adj_267), .C(n1061[22]), 
         .D(n2022[13]), .Z(n10_adj_269)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_160.init = 16'hfeee;
    LUT4 mux_220_Mux_22_i7_4_lut (.A(n67515), .B(\hidden_outputs[4] [22]), 
         .C(n[2]), .D(n70842), .Z(n3742[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_22_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_161 (.A(n3742[22]), .B(n10_adj_269), .C(n16_adj_268), 
         .D(n2022[35]), .Z(n63157)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_161.init = 16'hfefc;
    LUT4 mux_75_Mux_21_i7_4_lut (.A(n67299), .B(\temp_outputs[4] [21]), 
         .C(i[2]), .D(n17802), .Z(n1028[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_21_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i22_3_lut (.A(n1028[21]), .B(n1027[21]), .C(n70712), .Z(n1061[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i22_3_lut.init = 16'hacac;
    LUT4 select_455_Select_25_i32_2_lut (.A(sram_output_B[25]), .B(n2022[31]), 
         .Z(n32_adj_270)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_25_i32_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_162 (.A(f[21]), .B(n2448[21]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_271)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_162.init = 16'heca0;
    LUT4 select_460_Select_21_i16_2_lut (.A(e[21]), .B(n2022[15]), .Z(n16_adj_272)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_21_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_163 (.A(n17634), .B(n8_adj_271), .C(n1061[21]), 
         .D(n2022[13]), .Z(n10_adj_273)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_163.init = 16'hfeee;
    LUT4 mux_220_Mux_21_i7_4_lut (.A(n67512), .B(\hidden_outputs[4] [21]), 
         .C(n[2]), .D(n70842), .Z(n3742[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_21_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_164 (.A(n3742[21]), .B(n10_adj_273), .C(n16_adj_272), 
         .D(n2022[35]), .Z(n63161)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_164.init = 16'hfefc;
    LUT4 mux_75_Mux_20_i7_4_lut (.A(n67266), .B(\temp_outputs[4] [20]), 
         .C(i[2]), .D(n17802), .Z(n1028[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_20_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i21_3_lut (.A(n1028[20]), .B(n1027[20]), .C(n70712), .Z(n1061[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i21_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_165 (.A(f[20]), .B(n2448[20]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_274)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_165.init = 16'heca0;
    LUT4 i1_4_lut_adj_166 (.A(\mlp_outputs[1] [25]), .B(n70809), .C(float_alu_c[25]), 
         .D(o[0]), .Z(n23501)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_166.init = 16'hc088;
    LUT4 i2_4_lut_adj_167 (.A(n23501), .B(n32_adj_270), .C(\mlp_outputs[1] [25]), 
         .D(n2022[39]), .Z(n63240)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_167.init = 16'hfeee;
    LUT4 select_460_Select_20_i16_2_lut (.A(e[20]), .B(n2022[15]), .Z(n16_adj_275)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_20_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_168 (.A(n17619), .B(n8_adj_274), .C(n1061[20]), 
         .D(n2022[13]), .Z(n10_adj_276)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_168.init = 16'hfeee;
    LUT4 mux_220_Mux_20_i7_4_lut (.A(n67509), .B(\hidden_outputs[4] [20]), 
         .C(n[2]), .D(n70842), .Z(n3742[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_20_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_169 (.A(n3742[20]), .B(n10_adj_276), .C(n16_adj_275), 
         .D(n2022[35]), .Z(n63160)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_169.init = 16'hfefc;
    LUT4 mux_75_Mux_19_i7_4_lut (.A(n67302), .B(\temp_outputs[4] [19]), 
         .C(i[2]), .D(n17802), .Z(n1028[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_19_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i20_3_lut (.A(n1028[19]), .B(n1027[19]), .C(n70712), .Z(n1061[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i20_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_170 (.A(f[19]), .B(n2448[19]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_277)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_170.init = 16'heca0;
    LUT4 select_460_Select_19_i16_2_lut (.A(e[19]), .B(n2022[15]), .Z(n16_adj_278)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_19_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_171 (.A(n17405), .B(n8_adj_277), .C(n1061[19]), 
         .D(n2022[13]), .Z(n10_adj_279)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_171.init = 16'hfeee;
    LUT4 select_455_Select_26_i32_2_lut (.A(sram_output_B[26]), .B(n2022[31]), 
         .Z(n32_adj_280)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_26_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_172 (.A(\mlp_outputs[1] [26]), .B(n70809), .C(float_alu_c[26]), 
         .D(o[0]), .Z(n22808)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_172.init = 16'hc088;
    LUT4 i1_4_lut_adj_173 (.A(n32_adj_280), .B(n22808), .C(\mlp_outputs[1] [26]), 
         .D(n2022[39]), .Z(n66452)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_173.init = 16'hfeee;
    LUT4 select_455_Select_27_i32_2_lut (.A(sram_output_B[27]), .B(n2022[31]), 
         .Z(n32_adj_281)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_455_Select_27_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_174 (.A(\mlp_outputs[1] [27]), .B(n70809), .C(float_alu_c[27]), 
         .D(o[0]), .Z(n23498)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_174.init = 16'hc088;
    LUT4 mux_220_Mux_19_i7_4_lut (.A(n67506), .B(\hidden_outputs[4] [19]), 
         .C(n[2]), .D(n70842), .Z(n3742[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_19_i7_4_lut.init = 16'h0aca;
    LUT4 i2_4_lut_adj_175 (.A(n23498), .B(n32_adj_281), .C(\mlp_outputs[1] [27]), 
         .D(n2022[39]), .Z(n63239)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_175.init = 16'hfeee;
    LUT4 i5_4_lut_adj_176 (.A(n3742[19]), .B(n10_adj_279), .C(n16_adj_278), 
         .D(n2022[35]), .Z(n63245)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_176.init = 16'hfefc;
    LUT4 select_456_Select_28_i32_2_lut (.A(sram_output_B[28]), .B(n2022[31]), 
         .Z(n32_adj_282)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_28_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_177 (.A(\mlp_outputs[1] [28]), .B(n70809), .C(float_alu_c[28]), 
         .D(o[0]), .Z(n22868)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_177.init = 16'hc088;
    LUT4 i1_4_lut_adj_178 (.A(n32_adj_282), .B(n22868), .C(\mlp_outputs[1] [28]), 
         .D(n2022[39]), .Z(n66432)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_178.init = 16'hfeee;
    LUT4 select_456_Select_29_i32_2_lut (.A(sram_output_B[29]), .B(n2022[31]), 
         .Z(n32_adj_283)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_29_i32_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_179 (.A(\mlp_outputs[1] [29]), .B(n70809), .C(float_alu_c[29]), 
         .D(o[0]), .Z(n23414)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_179.init = 16'hc088;
    LUT4 i2_4_lut_adj_180 (.A(n23414), .B(n32_adj_283), .C(\mlp_outputs[1] [29]), 
         .D(n2022[39]), .Z(n63210)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_180.init = 16'hfeee;
    LUT4 mux_75_Mux_18_i7_4_lut (.A(n67305), .B(\temp_outputs[4] [18]), 
         .C(i[2]), .D(n17802), .Z(n1028[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_18_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i19_3_lut (.A(n1028[18]), .B(n1027[18]), .C(n70712), .Z(n1061[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i19_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_181 (.A(f[18]), .B(n2448[18]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_284)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_181.init = 16'heca0;
    PFUMX i54487 (.BLUT(n67396), .ALUT(n67397), .C0(h[1]), .Z(n67398));
    LUT4 select_456_Select_30_i32_2_lut (.A(sram_output_B[30]), .B(n2022[31]), 
         .Z(n32_adj_285)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_30_i32_2_lut.init = 16'h8888;
    LUT4 select_460_Select_18_i16_2_lut (.A(e[18]), .B(n2022[15]), .Z(n16_adj_286)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_18_i16_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_182 (.A(\mlp_outputs[1] [30]), .B(n70809), .C(float_alu_c[30]), 
         .D(o[0]), .Z(n23393)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_182.init = 16'hc088;
    LUT4 i1_4_lut_adj_183 (.A(n32_adj_285), .B(\mlp_outputs[1] [30]), .C(n23393), 
         .D(n2022[39]), .Z(n66376)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_183.init = 16'hfefa;
    LUT4 i4_4_lut_adj_184 (.A(n17365), .B(n8_adj_284), .C(n1061[18]), 
         .D(n2022[13]), .Z(n10_adj_287)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_184.init = 16'hfeee;
    LUT4 mux_220_Mux_18_i7_4_lut (.A(n67503), .B(\hidden_outputs[4] [18]), 
         .C(n[2]), .D(n70842), .Z(n3742[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_18_i7_4_lut.init = 16'h0aca;
    LUT4 select_456_Select_31_i32_2_lut (.A(sram_output_B[31]), .B(n2022[31]), 
         .Z(n32_adj_289)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_31_i32_2_lut.init = 16'h8888;
    LUT4 i20_2_lut (.A(o[0]), .B(\mlp_outputs[1] [31]), .Z(n10_adj_290)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i20_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_185 (.A(\mlp_outputs[1] [31]), .B(n70809), .C(float_alu_c[31]), 
         .D(o[0]), .Z(n23396)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_185.init = 16'hc088;
    LUT4 i2_4_lut_adj_186 (.A(n23396), .B(n32_adj_289), .C(n2022[39]), 
         .D(n10_adj_290), .Z(n63201)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_186.init = 16'hfeee;
    LUT4 i5_4_lut_adj_187 (.A(n3742[18]), .B(n10_adj_287), .C(n16_adj_286), 
         .D(n2022[35]), .Z(n63165)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_187.init = 16'hfefc;
    LUT4 mux_75_Mux_17_i7_4_lut (.A(n67308), .B(\temp_outputs[4] [17]), 
         .C(i[2]), .D(n17802), .Z(n1028[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_17_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i18_3_lut (.A(n1028[17]), .B(n1027[17]), .C(n70712), .Z(n1061[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i18_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_188 (.A(f[17]), .B(n2448[17]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_291)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_188.init = 16'heca0;
    FD1P3AX hidden_outputs_0__i0_i2 (.D(n66528), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [2]));
    defparam hidden_outputs_0__i0_i2.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i3 (.D(n66548), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [3]));
    defparam hidden_outputs_0__i0_i3.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i4 (.D(n63002), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [4]));
    defparam hidden_outputs_0__i0_i4.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i5 (.D(n66420), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [5]));
    defparam hidden_outputs_0__i0_i5.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i6 (.D(n66422), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [6]));
    defparam hidden_outputs_0__i0_i6.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i7 (.D(n63000), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [7]));
    defparam hidden_outputs_0__i0_i7.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i8 (.D(n66428), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [8]));
    defparam hidden_outputs_0__i0_i8.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i9 (.D(n66426), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [9]));
    defparam hidden_outputs_0__i0_i9.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i10 (.D(n62988), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [10]));
    defparam hidden_outputs_0__i0_i10.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i11 (.D(n63207), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [11]));
    defparam hidden_outputs_0__i0_i11.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i12 (.D(n66444), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [12]));
    defparam hidden_outputs_0__i0_i12.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i13 (.D(n63024), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [13]));
    defparam hidden_outputs_0__i0_i13.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i14 (.D(n63027), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [14]));
    defparam hidden_outputs_0__i0_i14.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i15 (.D(n66374), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [15]));
    defparam hidden_outputs_0__i0_i15.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i16 (.D(n62875), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [16]));
    defparam hidden_outputs_0__i0_i16.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i17 (.D(n63223), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [17]));
    defparam hidden_outputs_0__i0_i17.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i18 (.D(n63224), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [18]));
    defparam hidden_outputs_0__i0_i18.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i19 (.D(n63049), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [19]));
    defparam hidden_outputs_0__i0_i19.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i20 (.D(n66356), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [20]));
    defparam hidden_outputs_0__i0_i20.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i21 (.D(n62975), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [21]));
    defparam hidden_outputs_0__i0_i21.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i22 (.D(n66402), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [22]));
    defparam hidden_outputs_0__i0_i22.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i23 (.D(n66448), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [23]));
    defparam hidden_outputs_0__i0_i23.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i24 (.D(n63046), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [24]));
    defparam hidden_outputs_0__i0_i24.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i25 (.D(n62971), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [25]));
    defparam hidden_outputs_0__i0_i25.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i26 (.D(n66346), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [26]));
    defparam hidden_outputs_0__i0_i26.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i27 (.D(n66312), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [27]));
    defparam hidden_outputs_0__i0_i27.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i28 (.D(n63095), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [28]));
    defparam hidden_outputs_0__i0_i28.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i29 (.D(n63052), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [29]));
    defparam hidden_outputs_0__i0_i29.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i30 (.D(n66538), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [30]));
    defparam hidden_outputs_0__i0_i30.GSR = "DISABLED";
    FD1P3AX hidden_outputs_0__i0_i31 (.D(n63060), .SP(n23658), .CK(clock), 
            .Q(\hidden_outputs[0] [31]));
    defparam hidden_outputs_0__i0_i31.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i1 (.D(n66284), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [1]));
    defparam hidden_outputs_1__i0_i1.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i2 (.D(n62912), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [2]));
    defparam hidden_outputs_1__i0_i2.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i3 (.D(n66278), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [3]));
    defparam hidden_outputs_1__i0_i3.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i4 (.D(n66514), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [4]));
    defparam hidden_outputs_1__i0_i4.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i5 (.D(n63076), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [5]));
    defparam hidden_outputs_1__i0_i5.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i6 (.D(n62909), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [6]));
    defparam hidden_outputs_1__i0_i6.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i7 (.D(n66540), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [7]));
    defparam hidden_outputs_1__i0_i7.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i8 (.D(n66542), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [8]));
    defparam hidden_outputs_1__i0_i8.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i9 (.D(n62907), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [9]));
    defparam hidden_outputs_1__i0_i9.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i10 (.D(n62855), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [10]));
    defparam hidden_outputs_1__i0_i10.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i11 (.D(n66314), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [11]));
    defparam hidden_outputs_1__i0_i11.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i12 (.D(n66518), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [12]));
    defparam hidden_outputs_1__i0_i12.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i13 (.D(n66562), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [13]));
    defparam hidden_outputs_1__i0_i13.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i14 (.D(n62905), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [14]));
    defparam hidden_outputs_1__i0_i14.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i15 (.D(n66520), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [15]));
    defparam hidden_outputs_1__i0_i15.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i16 (.D(n66410), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [16]));
    defparam hidden_outputs_1__i0_i16.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i17 (.D(n66308), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [17]));
    defparam hidden_outputs_1__i0_i17.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i18 (.D(n66370), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [18]));
    defparam hidden_outputs_1__i0_i18.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i19 (.D(n66382), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [19]));
    defparam hidden_outputs_1__i0_i19.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i20 (.D(n63194), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [20]));
    defparam hidden_outputs_1__i0_i20.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i21 (.D(n66414), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [21]));
    defparam hidden_outputs_1__i0_i21.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i22 (.D(n66380), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [22]));
    defparam hidden_outputs_1__i0_i22.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i23 (.D(n66416), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [23]));
    defparam hidden_outputs_1__i0_i23.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i24 (.D(n63197), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [24]));
    defparam hidden_outputs_1__i0_i24.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i25 (.D(n63004), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [25]));
    defparam hidden_outputs_1__i0_i25.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i26 (.D(n66378), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [26]));
    defparam hidden_outputs_1__i0_i26.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i27 (.D(n66418), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [27]));
    defparam hidden_outputs_1__i0_i27.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i28 (.D(n66332), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [28]));
    defparam hidden_outputs_1__i0_i28.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i29 (.D(n62899), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [29]));
    defparam hidden_outputs_1__i0_i29.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i30 (.D(n66430), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [30]));
    defparam hidden_outputs_1__i0_i30.GSR = "DISABLED";
    FD1P3AX hidden_outputs_1__i0_i31 (.D(n66324), .SP(n23659), .CK(clock), 
            .Q(\hidden_outputs[1] [31]));
    defparam hidden_outputs_1__i0_i31.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i1 (.D(n66296), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [1]));
    defparam hidden_outputs_2__i0_i1.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i2 (.D(n62932), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [2]));
    defparam hidden_outputs_2__i0_i2.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i3 (.D(n66492), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [3]));
    defparam hidden_outputs_2__i0_i3.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i4 (.D(n63093), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [4]));
    defparam hidden_outputs_2__i0_i4.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i5 (.D(n66500), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [5]));
    defparam hidden_outputs_2__i0_i5.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i6 (.D(n63094), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [6]));
    defparam hidden_outputs_2__i0_i6.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i7 (.D(n62925), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [7]));
    defparam hidden_outputs_2__i0_i7.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i8 (.D(n66502), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [8]));
    defparam hidden_outputs_2__i0_i8.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i9 (.D(n66304), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [9]));
    defparam hidden_outputs_2__i0_i9.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i10 (.D(n63091), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [10]));
    defparam hidden_outputs_2__i0_i10.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i11 (.D(n66504), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [11]));
    defparam hidden_outputs_2__i0_i11.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i12 (.D(n66272), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [12]));
    defparam hidden_outputs_2__i0_i12.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i13 (.D(n62922), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [13]));
    defparam hidden_outputs_2__i0_i13.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i14 (.D(n66274), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [14]));
    defparam hidden_outputs_2__i0_i14.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i15 (.D(n63192), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [15]));
    defparam hidden_outputs_2__i0_i15.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i16 (.D(n66506), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [16]));
    defparam hidden_outputs_2__i0_i16.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i17 (.D(n63083), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [17]));
    defparam hidden_outputs_2__i0_i17.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i18 (.D(n62920), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [18]));
    defparam hidden_outputs_2__i0_i18.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i19 (.D(n66290), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [19]));
    defparam hidden_outputs_2__i0_i19.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i20 (.D(n66406), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [20]));
    defparam hidden_outputs_2__i0_i20.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i21 (.D(n63078), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [21]));
    defparam hidden_outputs_2__i0_i21.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i22 (.D(n66508), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [22]));
    defparam hidden_outputs_2__i0_i22.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i23 (.D(n66294), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [23]));
    defparam hidden_outputs_2__i0_i23.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i24 (.D(n62916), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [24]));
    defparam hidden_outputs_2__i0_i24.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i25 (.D(n63085), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [25]));
    defparam hidden_outputs_2__i0_i25.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i26 (.D(n66510), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [26]));
    defparam hidden_outputs_2__i0_i26.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i27 (.D(n66288), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [27]));
    defparam hidden_outputs_2__i0_i27.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i28 (.D(n66266), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [28]));
    defparam hidden_outputs_2__i0_i28.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i29 (.D(n62914), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [29]));
    defparam hidden_outputs_2__i0_i29.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i30 (.D(n63080), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [30]));
    defparam hidden_outputs_2__i0_i30.GSR = "DISABLED";
    FD1P3AX hidden_outputs_2__i0_i31 (.D(n66512), .SP(n23660), .CK(clock), 
            .Q(\hidden_outputs[2] [31]));
    defparam hidden_outputs_2__i0_i31.GSR = "DISABLED";
    LUT4 select_460_Select_17_i16_2_lut (.A(e[17]), .B(n2022[15]), .Z(n16_adj_292)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_17_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_189 (.A(n17345), .B(n8_adj_291), .C(n1061[17]), 
         .D(n2022[13]), .Z(n10_adj_293)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_189.init = 16'hfeee;
    LUT4 mux_220_Mux_17_i7_4_lut (.A(n67500), .B(\hidden_outputs[4] [17]), 
         .C(n[2]), .D(n70842), .Z(n3742[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_17_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_190 (.A(n3742[17]), .B(n10_adj_293), .C(n16_adj_292), 
         .D(n2022[35]), .Z(n63253)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_190.init = 16'hfefc;
    LUT4 mux_75_Mux_16_i7_4_lut (.A(n67311), .B(\temp_outputs[4] [16]), 
         .C(i[2]), .D(n17802), .Z(n1028[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_16_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i17_3_lut (.A(n1028[16]), .B(n1027[16]), .C(n70712), .Z(n1061[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i17_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_191 (.A(f[16]), .B(n2448[16]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_294)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_191.init = 16'heca0;
    PFUMX i54490 (.BLUT(n67399), .ALUT(n67400), .C0(h[1]), .Z(n67401));
    LUT4 select_460_Select_16_i16_2_lut (.A(e[16]), .B(n2022[15]), .Z(n16_adj_295)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_16_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_192 (.A(n17309), .B(n8_adj_294), .C(n1061[16]), 
         .D(n2022[13]), .Z(n10_adj_296)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_192.init = 16'hfeee;
    LUT4 mux_220_Mux_16_i7_4_lut (.A(n67497), .B(\hidden_outputs[4] [16]), 
         .C(n[2]), .D(n70842), .Z(n3742[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_16_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_193 (.A(n3742[16]), .B(n10_adj_296), .C(n16_adj_295), 
         .D(n2022[35]), .Z(n63153)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_193.init = 16'hfefc;
    LUT4 mux_75_Mux_15_i7_4_lut (.A(n67314), .B(\temp_outputs[4] [15]), 
         .C(i[2]), .D(n17802), .Z(n1028[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_15_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i16_3_lut (.A(n1028[15]), .B(n1027[15]), .C(n70712), .Z(n1061[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i16_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_194 (.A(f[15]), .B(n2448[15]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_297)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_194.init = 16'heca0;
    LUT4 select_460_Select_15_i16_2_lut (.A(e[15]), .B(n2022[15]), .Z(n16_adj_298)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_15_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_195 (.A(n17887), .B(n8_adj_297), .C(n1061[15]), 
         .D(n2022[13]), .Z(n10_adj_299)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_195.init = 16'hfeee;
    LUT4 mux_220_Mux_15_i7_4_lut (.A(n67494), .B(\hidden_outputs[4] [15]), 
         .C(n[2]), .D(n70842), .Z(n3742[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_15_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_196 (.A(n3742[15]), .B(n10_adj_299), .C(n16_adj_298), 
         .D(n2022[35]), .Z(n63146)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_196.init = 16'hfefc;
    LUT4 i1_4_lut_adj_197 (.A(n70822), .B(n2022[31]), .C(n2082), .D(n4_adj_72), 
         .Z(n46466)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_197.init = 16'h2220;
    LUT4 select_456_Select_0_i32_2_lut (.A(sram_output_B[0]), .B(n2022[31]), 
         .Z(n32_adj_111)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_456_Select_0_i32_2_lut.init = 16'h8888;
    LUT4 mux_75_Mux_14_i7_4_lut (.A(n67317), .B(\temp_outputs[4] [14]), 
         .C(i[2]), .D(n17802), .Z(n1028[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_14_i7_4_lut.init = 16'h0aca;
    LUT4 i4_4_lut_adj_198 (.A(n2022[43]), .B(n2022[47]), .C(n2022[49]), 
         .D(n2022[41]), .Z(n10_adj_71)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut_adj_198.init = 16'hfffe;
    LUT4 mux_76_i15_3_lut (.A(n1028[14]), .B(n1027[14]), .C(n70712), .Z(n1061[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i15_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_199 (.A(f[14]), .B(n2448[14]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_300)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_199.init = 16'heca0;
    FD1P3AX hidden_outputs_3__i0_i1 (.D(n66472), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [1]));
    defparam hidden_outputs_3__i0_i1.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i2 (.D(n66486), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [2]));
    defparam hidden_outputs_3__i0_i2.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i3 (.D(n62949), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [3]));
    defparam hidden_outputs_3__i0_i3.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i4 (.D(n62948), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [4]));
    defparam hidden_outputs_3__i0_i4.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i5 (.D(n66476), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [5]));
    defparam hidden_outputs_3__i0_i5.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i6 (.D(n63168), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [6]));
    defparam hidden_outputs_3__i0_i6.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i7 (.D(n62946), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [7]));
    defparam hidden_outputs_3__i0_i7.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i8 (.D(n66394), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [8]));
    defparam hidden_outputs_3__i0_i8.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i9 (.D(n66552), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [9]));
    defparam hidden_outputs_3__i0_i9.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i10 (.D(n66478), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [10]));
    defparam hidden_outputs_3__i0_i10.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i11 (.D(n66392), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [11]));
    defparam hidden_outputs_3__i0_i11.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i12 (.D(n62944), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [12]));
    defparam hidden_outputs_3__i0_i12.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i13 (.D(n63173), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [13]));
    defparam hidden_outputs_3__i0_i13.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i14 (.D(n66554), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [14]));
    defparam hidden_outputs_3__i0_i14.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i15 (.D(n66480), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [15]));
    defparam hidden_outputs_3__i0_i15.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i16 (.D(n63199), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [16]));
    defparam hidden_outputs_3__i0_i16.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i17 (.D(n62942), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [17]));
    defparam hidden_outputs_3__i0_i17.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i18 (.D(n66372), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [18]));
    defparam hidden_outputs_3__i0_i18.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i19 (.D(n66482), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [19]));
    defparam hidden_outputs_3__i0_i19.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i20 (.D(n66496), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [20]));
    defparam hidden_outputs_3__i0_i20.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i21 (.D(n62940), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [21]));
    defparam hidden_outputs_3__i0_i21.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i22 (.D(n66358), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [22]));
    defparam hidden_outputs_3__i0_i22.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i23 (.D(n62938), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [23]));
    defparam hidden_outputs_3__i0_i23.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i24 (.D(n66354), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [24]));
    defparam hidden_outputs_3__i0_i24.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i25 (.D(n62937), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [25]));
    defparam hidden_outputs_3__i0_i25.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i26 (.D(n66352), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [26]));
    defparam hidden_outputs_3__i0_i26.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i27 (.D(n66488), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [27]));
    defparam hidden_outputs_3__i0_i27.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i28 (.D(n66544), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [28]));
    defparam hidden_outputs_3__i0_i28.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i29 (.D(n62934), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [29]));
    defparam hidden_outputs_3__i0_i29.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i30 (.D(n63252), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [30]));
    defparam hidden_outputs_3__i0_i30.GSR = "DISABLED";
    FD1P3AX hidden_outputs_3__i0_i31 (.D(n66490), .SP(n23663), .CK(clock), 
            .Q(\hidden_outputs[3] [31]));
    defparam hidden_outputs_3__i0_i31.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i1 (.D(n63118), .SP(n23664), .CK(clock), .Q(float_alu_b[1]));
    defparam float_alu_b_i0_i1.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i2 (.D(n63117), .SP(n23664), .CK(clock), .Q(float_alu_b[2]));
    defparam float_alu_b_i0_i2.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i3 (.D(n63132), .SP(n23664), .CK(clock), .Q(float_alu_b[3]));
    defparam float_alu_b_i0_i3.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i4 (.D(n63134), .SP(n23664), .CK(clock), .Q(float_alu_b[4]));
    defparam float_alu_b_i0_i4.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i5 (.D(n63149), .SP(n23664), .CK(clock), .Q(float_alu_b[5]));
    defparam float_alu_b_i0_i5.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i6 (.D(n63256), .SP(n23664), .CK(clock), .Q(float_alu_b[6]));
    defparam float_alu_b_i0_i6.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i7 (.D(n63137), .SP(n23664), .CK(clock), .Q(float_alu_b[7]));
    defparam float_alu_b_i0_i7.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i8 (.D(n63136), .SP(n23664), .CK(clock), .Q(float_alu_b[8]));
    defparam float_alu_b_i0_i8.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i9 (.D(n63143), .SP(n23664), .CK(clock), .Q(float_alu_b[9]));
    defparam float_alu_b_i0_i9.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i10 (.D(n63140), .SP(n23664), .CK(clock), .Q(float_alu_b[10]));
    defparam float_alu_b_i0_i10.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i11 (.D(n63141), .SP(n23664), .CK(clock), .Q(float_alu_b[11]));
    defparam float_alu_b_i0_i11.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i12 (.D(n63144), .SP(n23664), .CK(clock), .Q(float_alu_b[12]));
    defparam float_alu_b_i0_i12.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i13 (.D(n63196), .SP(n23664), .CK(clock), .Q(float_alu_b[13]));
    defparam float_alu_b_i0_i13.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i14 (.D(n63145), .SP(n23664), .CK(clock), .Q(float_alu_b[14]));
    defparam float_alu_b_i0_i14.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i15 (.D(n63146), .SP(n23664), .CK(clock), .Q(float_alu_b[15]));
    defparam float_alu_b_i0_i15.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i16 (.D(n63153), .SP(n23664), .CK(clock), .Q(float_alu_b[16]));
    defparam float_alu_b_i0_i16.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i17 (.D(n63253), .SP(n23664), .CK(clock), .Q(float_alu_b[17]));
    defparam float_alu_b_i0_i17.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i18 (.D(n63165), .SP(n23664), .CK(clock), .Q(float_alu_b[18]));
    defparam float_alu_b_i0_i18.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i19 (.D(n63245), .SP(n23664), .CK(clock), .Q(float_alu_b[19]));
    defparam float_alu_b_i0_i19.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i20 (.D(n63160), .SP(n23664), .CK(clock), .Q(float_alu_b[20]));
    defparam float_alu_b_i0_i20.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i21 (.D(n63161), .SP(n23664), .CK(clock), .Q(float_alu_b[21]));
    defparam float_alu_b_i0_i21.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i22 (.D(n63157), .SP(n23664), .CK(clock), .Q(float_alu_b[22]));
    defparam float_alu_b_i0_i22.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i23 (.D(n63015), .SP(n23664), .CK(clock), .Q(float_alu_b[23]));
    defparam float_alu_b_i0_i23.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i25 (.D(n66404), .SP(n23664), .CK(clock), .Q(float_alu_b[25]));
    defparam float_alu_b_i0_i25.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i26 (.D(n66412), .SP(n23664), .CK(clock), .Q(float_alu_b[26]));
    defparam float_alu_b_i0_i26.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i27 (.D(n66310), .SP(n23664), .CK(clock), .Q(float_alu_b[27]));
    defparam float_alu_b_i0_i27.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i29 (.D(n66484), .SP(n23664), .CK(clock), .Q(float_alu_b[29]));
    defparam float_alu_b_i0_i29.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i30 (.D(n63151), .SP(n23664), .CK(clock), .Q(float_alu_b[30]));
    defparam float_alu_b_i0_i30.GSR = "DISABLED";
    FD1P3AX float_alu_b_i0_i31 (.D(n63021), .SP(n23664), .CK(clock), .Q(float_alu_b[31]));
    defparam float_alu_b_i0_i31.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i1 (.D(n66282), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [1]));
    defparam hidden_outputs_4__i0_i1.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i2 (.D(n66470), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [2]));
    defparam hidden_outputs_4__i0_i2.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i3 (.D(n66344), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [3]));
    defparam hidden_outputs_4__i0_i3.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i4 (.D(n66516), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [4]));
    defparam hidden_outputs_4__i0_i4.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i5 (.D(n62864), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [5]));
    defparam hidden_outputs_4__i0_i5.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i6 (.D(n66546), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [6]));
    defparam hidden_outputs_4__i0_i6.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i7 (.D(n66328), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [7]));
    defparam hidden_outputs_4__i0_i7.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i8 (.D(n66550), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [8]));
    defparam hidden_outputs_4__i0_i8.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i9 (.D(n66424), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [9]));
    defparam hidden_outputs_4__i0_i9.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i10 (.D(n66286), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [10]));
    defparam hidden_outputs_4__i0_i10.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i11 (.D(n66450), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [11]));
    defparam hidden_outputs_4__i0_i11.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i12 (.D(n66268), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [12]));
    defparam hidden_outputs_4__i0_i12.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i13 (.D(n66462), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [13]));
    defparam hidden_outputs_4__i0_i13.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i14 (.D(n66536), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [14]));
    defparam hidden_outputs_4__i0_i14.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i15 (.D(n66276), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [15]));
    defparam hidden_outputs_4__i0_i15.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i16 (.D(n66398), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [16]));
    defparam hidden_outputs_4__i0_i16.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i17 (.D(n66330), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [17]));
    defparam hidden_outputs_4__i0_i17.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i18 (.D(n66388), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [18]));
    defparam hidden_outputs_4__i0_i18.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i19 (.D(n66270), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [19]));
    defparam hidden_outputs_4__i0_i19.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i20 (.D(n66302), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [20]));
    defparam hidden_outputs_4__i0_i20.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i21 (.D(n66318), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [21]));
    defparam hidden_outputs_4__i0_i21.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i22 (.D(n63014), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [22]));
    defparam hidden_outputs_4__i0_i22.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i23 (.D(n63190), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [23]));
    defparam hidden_outputs_4__i0_i23.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i24 (.D(n66360), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [24]));
    defparam hidden_outputs_4__i0_i24.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i25 (.D(n66498), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [25]));
    defparam hidden_outputs_4__i0_i25.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i26 (.D(n66326), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [26]));
    defparam hidden_outputs_4__i0_i26.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i27 (.D(n66408), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [27]));
    defparam hidden_outputs_4__i0_i27.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i28 (.D(n62953), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [28]));
    defparam hidden_outputs_4__i0_i28.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i29 (.D(n66384), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [29]));
    defparam hidden_outputs_4__i0_i29.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i30 (.D(n63065), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [30]));
    defparam hidden_outputs_4__i0_i30.GSR = "DISABLED";
    FD1P3AX hidden_outputs_4__i0_i31 (.D(n62951), .SP(n23665), .CK(clock), 
            .Q(\hidden_outputs[4] [31]));
    defparam hidden_outputs_4__i0_i31.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_200 (.A(\mlp_outputs[0] [0]), .B(n70809), .C(float_alu_c[0]), 
         .D(o[0]), .Z(n23357)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_200.init = 16'h88c0;
    PFUMX i54493 (.BLUT(n67402), .ALUT(n67403), .C0(h[1]), .Z(n67404));
    LUT4 i1_4_lut_adj_201 (.A(n32_adj_111), .B(\mlp_outputs[0] [0]), .C(n23357), 
         .D(n2022[39]), .Z(n66280)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_201.init = 16'hfefa;
    LUT4 select_460_Select_14_i16_2_lut (.A(e[14]), .B(n2022[15]), .Z(n16_adj_301)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_14_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_202 (.A(n17567), .B(n8_adj_300), .C(n1061[14]), 
         .D(n2022[13]), .Z(n10_adj_302)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_202.init = 16'hfeee;
    LUT4 mux_220_Mux_14_i7_4_lut (.A(n67491), .B(\hidden_outputs[4] [14]), 
         .C(n[2]), .D(n70842), .Z(n3742[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_14_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_203 (.A(n3742[14]), .B(n10_adj_302), .C(n16_adj_301), 
         .D(n2022[35]), .Z(n63145)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_203.init = 16'hfefc;
    PFUMX i54496 (.BLUT(n67405), .ALUT(n67406), .C0(h[1]), .Z(n67407));
    LUT4 mux_75_Mux_13_i7_4_lut (.A(n67320), .B(\temp_outputs[4] [13]), 
         .C(i[2]), .D(n17802), .Z(n1028[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_13_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i14_3_lut (.A(n1028[13]), .B(n1027[13]), .C(n70712), .Z(n1061[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i14_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_204 (.A(f[13]), .B(n2448[13]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_303)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_204.init = 16'heca0;
    LUT4 mux_141_Mux_0_i7_4_lut (.A(n67257), .B(\hidden_outputs[4] [0]), 
         .C(h[2]), .D(n70861), .Z(n2448[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_0_i7_4_lut.init = 16'h0aca;
    LUT4 select_460_Select_13_i16_2_lut (.A(e[13]), .B(n2022[15]), .Z(n16_adj_304)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_13_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_205 (.A(n17891), .B(n8_adj_303), .C(n1061[13]), 
         .D(n2022[13]), .Z(n10_adj_305)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_205.init = 16'hfeee;
    LUT4 mux_220_Mux_13_i7_4_lut (.A(n67488), .B(\hidden_outputs[4] [13]), 
         .C(n[2]), .D(n70842), .Z(n3742[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_13_i7_4_lut.init = 16'h0aca;
    PFUMX i54499 (.BLUT(n67408), .ALUT(n67409), .C0(h[1]), .Z(n67410));
    LUT4 i5_4_lut_adj_206 (.A(n3742[13]), .B(n10_adj_305), .C(n16_adj_304), 
         .D(n2022[35]), .Z(n63196)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_206.init = 16'hfefc;
    LUT4 i12324_2_lut_4_lut (.A(n70822), .B(n70859), .C(n70725), .D(n22276), 
         .Z(n24013)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;
    defparam i12324_2_lut_4_lut.init = 16'ha800;
    LUT4 mux_75_Mux_12_i7_4_lut (.A(n67323), .B(\temp_outputs[4] [12]), 
         .C(i[2]), .D(n17802), .Z(n1028[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_12_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i13_3_lut (.A(n1028[12]), .B(n1027[12]), .C(n70712), .Z(n1061[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i13_3_lut.init = 16'hacac;
    LUT4 mux_237_Mux_0_i1_3_lut (.A(\mlp_outputs[0] [0]), .B(\mlp_outputs[1] [0]), 
         .C(o[0]), .Z(n4478[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_0_i1_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_207 (.A(f[12]), .B(n2448[12]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_306)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_207.init = 16'heca0;
    LUT4 select_460_Select_12_i16_2_lut (.A(e[12]), .B(n2022[15]), .Z(n16_adj_307)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_12_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_208 (.A(n17895), .B(n8_adj_306), .C(n1061[12]), 
         .D(n2022[13]), .Z(n10_adj_308)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_208.init = 16'hfeee;
    LUT4 mux_220_Mux_12_i7_4_lut (.A(n67485), .B(\hidden_outputs[4] [12]), 
         .C(n[2]), .D(n70842), .Z(n3742[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_12_i7_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_adj_209 (.A(n2448[0]), .B(n23104), .Z(n22607)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_209.init = 16'h8888;
    LUT4 i5_4_lut_adj_210 (.A(n3742[12]), .B(n10_adj_308), .C(n16_adj_307), 
         .D(n2022[35]), .Z(n63144)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_210.init = 16'hfefc;
    LUT4 i2_4_lut_adj_211 (.A(n22607), .B(n22610), .C(weight[0]), .D(n70860), 
         .Z(n62900)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_211.init = 16'hfeee;
    LUT4 mux_75_Mux_11_i7_4_lut (.A(n67326), .B(\temp_outputs[4] [11]), 
         .C(i[2]), .D(n17802), .Z(n1028[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_11_i7_4_lut.init = 16'h0aca;
    PFUMX i54502 (.BLUT(n67411), .ALUT(n67412), .C0(h[1]), .Z(n67413));
    PFUMX i54505 (.BLUT(n67414), .ALUT(n67415), .C0(h[1]), .Z(n67416));
    LUT4 mux_76_i12_3_lut (.A(n1028[11]), .B(n1027[11]), .C(n70712), .Z(n1061[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i12_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_212 (.A(f[11]), .B(n2448[11]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_309)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_212.init = 16'heca0;
    LUT4 select_460_Select_11_i16_2_lut (.A(e[11]), .B(n2022[15]), .Z(n16_adj_310)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_11_i16_2_lut.init = 16'h8888;
    PFUMX i54508 (.BLUT(n67417), .ALUT(n67418), .C0(h[1]), .Z(n67419));
    PFUMX i54511 (.BLUT(n67420), .ALUT(n67421), .C0(h[1]), .Z(n67422));
    LUT4 i4_4_lut_adj_213 (.A(n17899), .B(n8_adj_309), .C(n1061[11]), 
         .D(n2022[13]), .Z(n10_adj_311)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_213.init = 16'hfeee;
    LUT4 mux_220_Mux_11_i7_4_lut (.A(n67482), .B(\hidden_outputs[4] [11]), 
         .C(n[2]), .D(n70842), .Z(n3742[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_11_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_214 (.A(n3742[11]), .B(n10_adj_311), .C(n16_adj_310), 
         .D(n2022[35]), .Z(n63141)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_214.init = 16'hfefc;
    LUT4 i7_2_lut (.A(o[2]), .B(o[29]), .Z(n39)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut.init = 16'heeee;
    LUT4 i19_4_lut_adj_215 (.A(o[19]), .B(o[8]), .C(o[20]), .D(o[12]), 
         .Z(n51)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_215.init = 16'hfffe;
    LUT4 i14_2_lut (.A(o[7]), .B(o[15]), .Z(n46)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut.init = 16'heeee;
    LUT4 i93_3_lut_4_lut (.A(n70723), .B(numL[31]), .C(n2022[28]), .D(n70724), 
         .Z(n2272)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i93_3_lut_4_lut.init = 16'hff20;
    LUT4 mux_75_Mux_10_i7_4_lut (.A(n67329), .B(\temp_outputs[4] [10]), 
         .C(i[2]), .D(n17802), .Z(n1028[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_10_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i11_3_lut (.A(n1028[10]), .B(n1027[10]), .C(n70712), .Z(n1061[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i11_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_216 (.A(f[10]), .B(n2448[10]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_312)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_216.init = 16'heca0;
    LUT4 i24_4_lut (.A(o[26]), .B(o[18]), .C(o[14]), .D(o[16]), .Z(n56_adj_313)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 select_460_Select_10_i16_2_lut (.A(e[10]), .B(n2022[15]), .Z(n16_adj_314)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_10_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_217 (.A(n17901), .B(n8_adj_312), .C(n1061[10]), 
         .D(n2022[13]), .Z(n10_adj_315)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_217.init = 16'hfeee;
    LUT4 mux_220_Mux_10_i7_4_lut (.A(n67479), .B(\hidden_outputs[4] [10]), 
         .C(n[2]), .D(n70842), .Z(n3742[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_10_i7_4_lut.init = 16'h0aca;
    LUT4 i10_2_lut (.A(o[30]), .B(o[25]), .Z(n42_adj_316)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i22_4_lut_adj_218 (.A(o[3]), .B(o[22]), .C(o[31]), .D(o[6]), 
         .Z(n1)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut_adj_218.init = 16'hfffe;
    LUT4 i5_4_lut_adj_219 (.A(n3742[10]), .B(n10_adj_315), .C(n16_adj_314), 
         .D(n2022[35]), .Z(n63140)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_219.init = 16'hfefc;
    LUT4 i28_4_lut (.A(o[9]), .B(n56_adj_313), .C(n46), .D(o[23]), .Z(n60_adj_317)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut.init = 16'hfffe;
    LUT4 i27929_2_lut_4_lut (.A(numL[0]), .B(n70723), .C(numL[31]), .D(n932), 
         .Z(n13947[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i27929_2_lut_4_lut.init = 16'hfe00;
    LUT4 i9_2_lut_adj_220 (.A(o[4]), .B(o[27]), .Z(n41)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut_adj_220.init = 16'heeee;
    LUT4 mux_75_Mux_9_i7_4_lut (.A(n67332), .B(\temp_outputs[4] [9]), .C(i[2]), 
         .D(n17802), .Z(n1028[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_9_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i10_3_lut (.A(n1028[9]), .B(n1027[9]), .C(n70712), .Z(n1061[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i10_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_221 (.A(f[9]), .B(n2448[9]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_318)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_221.init = 16'heca0;
    LUT4 i18_4_lut (.A(o[24]), .B(o[11]), .C(o[5]), .D(o[28]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i26_4_lut (.A(n51), .B(n39), .C(o[21]), .D(o[0]), .Z(n58_adj_319)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i26_4_lut.init = 16'hfeff;
    LUT4 i30_4_lut (.A(n41), .B(n60_adj_317), .C(n1), .D(n42_adj_316), 
         .Z(n62_adj_320)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut_adj_222 (.A(o[1]), .B(o[10]), .C(o[13]), .D(o[17]), 
         .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_222.init = 16'hfffe;
    LUT4 i31_4_lut (.A(n49), .B(n62_adj_320), .C(n58_adj_319), .D(n50), 
         .Z(n27496)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut.init = 16'hfffe;
    LUT4 select_460_Select_9_i16_2_lut (.A(e[9]), .B(n2022[15]), .Z(n16_adj_321)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_9_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_223 (.A(n17905), .B(n8_adj_318), .C(n1061[9]), .D(n2022[13]), 
         .Z(n10_adj_322)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_223.init = 16'hfeee;
    LUT4 mux_220_Mux_9_i7_4_lut (.A(n67476), .B(\hidden_outputs[4] [9]), 
         .C(n[2]), .D(n70842), .Z(n3742[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_9_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_224 (.A(n3742[9]), .B(n10_adj_322), .C(n16_adj_321), 
         .D(n2022[35]), .Z(n63143)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_224.init = 16'hfefc;
    LUT4 i29106_2_lut_4_lut (.A(numL[0]), .B(n70723), .C(numL[31]), .D(n930), 
         .Z(n13947[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i29106_2_lut_4_lut.init = 16'hfe00;
    LUT4 i29052_2_lut_4_lut (.A(numL[0]), .B(n70723), .C(numL[31]), .D(n236[3]), 
         .Z(n15041[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i29052_2_lut_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_adj_225 (.A(n2022[27]), .B(n2664), .Z(n2269)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_225.init = 16'h8888;
    LUT4 mux_75_Mux_8_i7_4_lut (.A(n67335), .B(\temp_outputs[4] [8]), .C(i[2]), 
         .D(n17802), .Z(n1028[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_8_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i9_3_lut (.A(n1028[8]), .B(n1027[8]), .C(n70712), .Z(n1061[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i9_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_226 (.A(f[8]), .B(n2448[8]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_323)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_226.init = 16'heca0;
    PFUMX i54514 (.BLUT(n67423), .ALUT(n67424), .C0(h[1]), .Z(n67425));
    LUT4 select_460_Select_8_i16_2_lut (.A(e[8]), .B(n2022[15]), .Z(n16_adj_324)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_8_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_227 (.A(n17909), .B(n8_adj_323), .C(n1061[8]), .D(n2022[13]), 
         .Z(n10_adj_325)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_227.init = 16'hfeee;
    LUT4 mux_220_Mux_8_i7_4_lut (.A(n67473), .B(\hidden_outputs[4] [8]), 
         .C(n[2]), .D(n70842), .Z(n3742[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_8_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_228 (.A(n3742[8]), .B(n10_adj_325), .C(n16_adj_324), 
         .D(n2022[35]), .Z(n63136)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_228.init = 16'hfefc;
    LUT4 mux_75_Mux_7_i7_4_lut (.A(n67338), .B(\temp_outputs[4] [7]), .C(i[2]), 
         .D(n17802), .Z(n1028[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_7_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i8_3_lut (.A(n1028[7]), .B(n1027[7]), .C(n70712), .Z(n1061[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i8_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_229 (.A(f[7]), .B(n2448[7]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_326)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_229.init = 16'heca0;
    LUT4 select_460_Select_7_i16_2_lut (.A(e[7]), .B(n2022[15]), .Z(n16_adj_327)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_7_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_230 (.A(n17911), .B(n8_adj_326), .C(n1061[7]), .D(n2022[13]), 
         .Z(n10_adj_328)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_230.init = 16'hfeee;
    LUT4 mux_220_Mux_7_i7_4_lut (.A(n67470), .B(\hidden_outputs[4] [7]), 
         .C(n[2]), .D(n70842), .Z(n3742[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_7_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_231 (.A(n3742[7]), .B(n10_adj_328), .C(n16_adj_327), 
         .D(n2022[35]), .Z(n63137)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_231.init = 16'hfefc;
    FD1P3IX addr_4653__i0 (.D(n134_adj_408[0]), .SP(n70769), .CD(n24023), 
            .CK(clock), .Q(addr[0]));
    defparam addr_4653__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut_adj_232 (.A(n236[0]), .B(n236[1]), .C(n70712), 
         .D(n236[2]), .Z(n66247)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_232.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_233 (.A(n236[0]), .B(n236[1]), .C(n70712), 
         .D(n236[2]), .Z(n65435)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_233.init = 16'hf080;
    LUT4 mux_75_Mux_6_i7_4_lut (.A(n67341), .B(\temp_outputs[4] [6]), .C(i[2]), 
         .D(n17802), .Z(n1028[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_6_i7_4_lut.init = 16'h0aca;
    LUT4 i2_3_lut_rep_738 (.A(n236[0]), .B(n236[1]), .C(n70712), .Z(n70708)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_738.init = 16'h8080;
    LUT4 mux_76_i7_3_lut (.A(n1028[6]), .B(n1027[6]), .C(n70712), .Z(n1061[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i7_3_lut.init = 16'hacac;
    LUT4 mux_141_Mux_29_i7_4_lut (.A(n67443), .B(\hidden_outputs[4] [29]), 
         .C(h[2]), .D(n70861), .Z(n2448[29])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_29_i7_4_lut.init = 16'h0aca;
    LUT4 i2_4_lut_adj_234 (.A(f[6]), .B(n2448[6]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_330)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_234.init = 16'heca0;
    LUT4 mux_237_Mux_29_i1_3_lut (.A(\mlp_outputs[0] [29]), .B(\mlp_outputs[1] [29]), 
         .C(o[0]), .Z(n4478[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_29_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_235 (.A(n23104), .B(n2448[29]), .Z(n23525)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_235.init = 16'h8888;
    LUT4 select_460_Select_6_i16_2_lut (.A(e[6]), .B(n2022[15]), .Z(n16_adj_331)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_6_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_236 (.A(n17881), .B(n8_adj_330), .C(n1061[6]), .D(n2022[13]), 
         .Z(n10_adj_332)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_236.init = 16'hfeee;
    LUT4 mux_220_Mux_6_i7_4_lut (.A(n67467), .B(\hidden_outputs[4] [6]), 
         .C(n[2]), .D(n70842), .Z(n3742[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_6_i7_4_lut.init = 16'h0aca;
    LUT4 i2_4_lut_adj_237 (.A(n23525), .B(n23528), .C(weight[29]), .D(n70860), 
         .Z(n63130)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_237.init = 16'hfeee;
    LUT4 i5_4_lut_adj_238 (.A(n3742[6]), .B(n10_adj_332), .C(n16_adj_331), 
         .D(n2022[35]), .Z(n63256)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_238.init = 16'hfefc;
    FD1S3AX No_Name_i2 (.D(\buf_x[84] ), .CK(clock), .Q(\buf_r[84] ));
    defparam No_Name_i2.GSR = "DISABLED";
    FD1S3AX No_Name_i3 (.D(\buf_x[85] ), .CK(clock), .Q(\buf_r[85] ));
    defparam No_Name_i3.GSR = "DISABLED";
    FD1S3AX No_Name_i4 (.D(\buf_x[86] ), .CK(clock), .Q(\buf_r[86] ));
    defparam No_Name_i4.GSR = "DISABLED";
    FD1S3AX No_Name_i5 (.D(\buf_x[87] ), .CK(clock), .Q(\buf_r[87] ));
    defparam No_Name_i5.GSR = "DISABLED";
    FD1S3AX No_Name_i6 (.D(\buf_x[88] ), .CK(clock), .Q(\buf_r[88] ));
    defparam No_Name_i6.GSR = "DISABLED";
    FD1S3AX No_Name_i7 (.D(\buf_x[89] ), .CK(clock), .Q(\buf_r[89] ));
    defparam No_Name_i7.GSR = "DISABLED";
    LUT4 mux_75_Mux_5_i7_4_lut (.A(n67344), .B(\temp_outputs[4] [5]), .C(i[2]), 
         .D(n17802), .Z(n1028[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_5_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i6_3_lut (.A(n1028[5]), .B(n1027[5]), .C(n70712), .Z(n1061[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i6_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_239 (.A(f[5]), .B(n2448[5]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_333)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_239.init = 16'heca0;
    LUT4 select_460_Select_5_i16_2_lut (.A(e[5]), .B(n2022[15]), .Z(n16_adj_334)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_5_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_240 (.A(n17919), .B(n8_adj_333), .C(n1061[5]), .D(n2022[13]), 
         .Z(n10_adj_335)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_240.init = 16'hfeee;
    LUT4 mux_220_Mux_5_i7_4_lut (.A(n67464), .B(\hidden_outputs[4] [5]), 
         .C(n[2]), .D(n70842), .Z(n3742[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_5_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_241 (.A(n3742[5]), .B(n10_adj_335), .C(n16_adj_334), 
         .D(n2022[35]), .Z(n63149)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_241.init = 16'hfefc;
    LUT4 mux_75_Mux_4_i7_4_lut (.A(n67347), .B(\temp_outputs[4] [4]), .C(i[2]), 
         .D(n17802), .Z(n1028[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_4_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i5_3_lut (.A(n1028[4]), .B(n1027[4]), .C(n70712), .Z(n1061[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i5_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_242 (.A(f[4]), .B(n2448[4]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_336)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_242.init = 16'heca0;
    LUT4 select_460_Select_4_i16_2_lut (.A(e[4]), .B(n2022[15]), .Z(n16_adj_337)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_4_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_243 (.A(n17921), .B(n8_adj_336), .C(n1061[4]), .D(n2022[13]), 
         .Z(n10_adj_338)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_243.init = 16'hfeee;
    LUT4 mux_220_Mux_4_i7_4_lut (.A(n67461), .B(\hidden_outputs[4] [4]), 
         .C(n[2]), .D(n70842), .Z(n3742[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_4_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_244 (.A(n3742[4]), .B(n10_adj_338), .C(n16_adj_337), 
         .D(n2022[35]), .Z(n63134)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_244.init = 16'hfefc;
    LUT4 i53913_3_lut_4_lut (.A(n236[2]), .B(n70708), .C(n236[3]), .D(n70712), 
         .Z(n66817)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C (D))))) */ ;
    defparam i53913_3_lut_4_lut.init = 16'h1e00;
    LUT4 mux_75_Mux_3_i7_4_lut (.A(n67350), .B(\temp_outputs[4] [3]), .C(i[2]), 
         .D(n17802), .Z(n1028[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_3_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i4_3_lut (.A(n1028[3]), .B(n1027[3]), .C(n70712), .Z(n1061[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i4_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_245 (.A(f[3]), .B(n2448[3]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_339)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_245.init = 16'heca0;
    LUT4 select_460_Select_3_i16_2_lut (.A(e[3]), .B(n2022[15]), .Z(n16_adj_340)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_3_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_246 (.A(n17925), .B(n8_adj_339), .C(n1061[3]), .D(n2022[13]), 
         .Z(n10_adj_341)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_246.init = 16'hfeee;
    LUT4 mux_220_Mux_3_i7_4_lut (.A(n67458), .B(\hidden_outputs[4] [3]), 
         .C(n[2]), .D(n70842), .Z(n3742[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_3_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_247 (.A(n3742[3]), .B(n10_adj_341), .C(n16_adj_340), 
         .D(n2022[35]), .Z(n63132)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_247.init = 16'hfefc;
    LUT4 mux_75_Mux_2_i7_4_lut (.A(n67353), .B(\temp_outputs[4] [2]), .C(i[2]), 
         .D(n17802), .Z(n1028[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_2_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i3_3_lut (.A(n1028[2]), .B(n1027[2]), .C(n70712), .Z(n1061[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i3_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_248 (.A(f[2]), .B(n2448[2]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_342)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_248.init = 16'heca0;
    LUT4 select_460_Select_2_i16_2_lut (.A(e[2]), .B(n2022[15]), .Z(n16_adj_343)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_2_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_249 (.A(n18121), .B(n8_adj_342), .C(n1061[2]), .D(n2022[13]), 
         .Z(n10_adj_344)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_249.init = 16'hfeee;
    LUT4 i1_2_lut_adj_250 (.A(n2022[22]), .B(n2022[44]), .Z(n22276)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_250.init = 16'heeee;
    LUT4 mux_220_Mux_2_i7_4_lut (.A(n67455), .B(\hidden_outputs[4] [2]), 
         .C(n[2]), .D(n70842), .Z(n3742[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_2_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_251 (.A(n3742[2]), .B(n10_adj_344), .C(n16_adj_343), 
         .D(n2022[35]), .Z(n63117)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_251.init = 16'hfefc;
    LUT4 i1_2_lut_adj_252 (.A(n2022[24]), .B(n2022[15]), .Z(n128)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_252.init = 16'heeee;
    LUT4 i3_4_lut_adj_253 (.A(n128), .B(n2022[26]), .C(n2022[18]), .D(n2022[20]), 
         .Z(n23104)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_253.init = 16'hfffe;
    LUT4 mux_141_Mux_28_i7_4_lut (.A(n67440), .B(\hidden_outputs[4] [28]), 
         .C(h[2]), .D(n70861), .Z(n2448[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_28_i7_4_lut.init = 16'h0aca;
    LUT4 mux_75_Mux_1_i7_4_lut (.A(n67356), .B(\temp_outputs[4] [1]), .C(i[2]), 
         .D(n17802), .Z(n1028[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_1_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i2_3_lut (.A(n1028[1]), .B(n1027[1]), .C(n70712), .Z(n1061[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i2_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_254 (.A(f[1]), .B(n2448[1]), .C(n2022[37]), .D(n17400), 
         .Z(n8_adj_345)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_254.init = 16'heca0;
    LUT4 i1_4_lut_rep_731 (.A(n2022[16]), .B(n23), .C(n1423), .D(n70712), 
         .Z(n70701)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i1_4_lut_rep_731.init = 16'ha022;
    LUT4 select_460_Select_1_i16_2_lut (.A(e[1]), .B(n2022[15]), .Z(n16_adj_346)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_1_i16_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_255 (.A(n18119), .B(n8_adj_345), .C(n1061[1]), .D(n2022[13]), 
         .Z(n10_adj_347)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_255.init = 16'hfeee;
    LUT4 mux_220_Mux_1_i7_4_lut (.A(n67452), .B(\hidden_outputs[4] [1]), 
         .C(n[2]), .D(n70842), .Z(n3742[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_1_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_28_i1_3_lut (.A(\mlp_outputs[0] [28]), .B(\mlp_outputs[1] [28]), 
         .C(o[0]), .Z(n4478[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_28_i1_3_lut.init = 16'hcaca;
    LUT4 i5_4_lut_adj_256 (.A(n3742[1]), .B(n10_adj_347), .C(n16_adj_346), 
         .D(n2022[35]), .Z(n63118)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_256.init = 16'hfefc;
    LUT4 i1_4_lut_rep_730 (.A(n2022[16]), .B(n23), .C(n1423), .D(n70712), 
         .Z(n70700)) /* synthesis lut_function=(!((B (C (D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_rep_730.init = 16'h0a88;
    LUT4 i1_2_lut_adj_257 (.A(n2448[28]), .B(n23104), .Z(n23345)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_257.init = 16'h8888;
    LUT4 i2_4_lut_adj_258 (.A(n23345), .B(n23348), .C(weight[28]), .D(n70860), 
         .Z(n63113)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_258.init = 16'hfeee;
    LUT4 i1_4_lut_adj_259 (.A(\hidden_outputs[3] [31]), .B(n22568), .C(float_alu_c[31]), 
         .D(n70785), .Z(n22682)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_259.init = 16'hc088;
    LUT4 i1_4_lut_adj_260 (.A(n10_adj_182), .B(n22682), .C(n1583), .D(n2022[17]), 
         .Z(n66490)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_260.init = 16'hfeee;
    LUT4 i1_4_lut_adj_261 (.A(\hidden_outputs[3] [30]), .B(n22568), .C(float_alu_c[30]), 
         .D(n70785), .Z(n23189)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_261.init = 16'hc088;
    LUT4 i2_4_lut_adj_262 (.A(n23189), .B(n10_adj_183), .C(\hidden_outputs[3] [30]), 
         .D(n2022[17]), .Z(n63252)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_262.init = 16'hfeee;
    LUT4 i1_4_lut_adj_263 (.A(\hidden_outputs[3] [29]), .B(n22568), .C(float_alu_c[29]), 
         .D(n70785), .Z(n22685)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_263.init = 16'hc088;
    LUT4 i2_4_lut_adj_264 (.A(n10_adj_185), .B(n22685), .C(\hidden_outputs[3] [29]), 
         .D(n2022[17]), .Z(n62934)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_264.init = 16'hfeee;
    LUT4 i1_4_lut_adj_265 (.A(\hidden_outputs[3] [28]), .B(n22568), .C(float_alu_c[28]), 
         .D(n70785), .Z(n23534)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_265.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_adj_266 (.A(n2022[38]), .B(n3922), .C(n2022[31]), 
         .Z(n2277)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_266.init = 16'hf2f2;
    LUT4 i1_4_lut_adj_267 (.A(n10_adj_186), .B(\hidden_outputs[3] [28]), 
         .C(n23534), .D(n2022[17]), .Z(n66544)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_267.init = 16'hfefa;
    LUT4 i1_4_lut_adj_268 (.A(\hidden_outputs[3] [27]), .B(n22568), .C(float_alu_c[27]), 
         .D(n70785), .Z(n22688)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_268.init = 16'hc088;
    PFUMX i54517 (.BLUT(n67426), .ALUT(n67427), .C0(h[1]), .Z(n67428));
    LUT4 i1_4_lut_adj_269 (.A(n10_adj_187), .B(n22688), .C(\hidden_outputs[3] [27]), 
         .D(n2022[17]), .Z(n66488)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_269.init = 16'hfeee;
    LUT4 i1_4_lut_rep_727_4_lut (.A(n2022[38]), .B(n3922), .C(n70822), 
         .D(n2022[31]), .Z(n70697)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C (D)))) */ ;
    defparam i1_4_lut_rep_727_4_lut.init = 16'h7020;
    LUT4 i1_4_lut_adj_270 (.A(\hidden_outputs[3] [26]), .B(n22568), .C(float_alu_c[26]), 
         .D(n70785), .Z(n23495)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_270.init = 16'hc088;
    LUT4 i1_4_lut_adj_271 (.A(n10_adj_188), .B(\hidden_outputs[3] [26]), 
         .C(n23495), .D(n2022[17]), .Z(n66352)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_271.init = 16'hfefa;
    LUT4 i1_4_lut_adj_272 (.A(\hidden_outputs[3] [25]), .B(n22568), .C(float_alu_c[25]), 
         .D(n70785), .Z(n22691)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_272.init = 16'hc088;
    LUT4 i2_4_lut_adj_273 (.A(n10_adj_189), .B(n22691), .C(\hidden_outputs[3] [25]), 
         .D(n2022[17]), .Z(n62937)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_273.init = 16'hfeee;
    LUT4 i1_4_lut_adj_274 (.A(\hidden_outputs[3] [24]), .B(n22568), .C(float_alu_c[24]), 
         .D(n70785), .Z(n23465)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_274.init = 16'hc088;
    LUT4 i1_4_lut_adj_275 (.A(n10_adj_190), .B(\hidden_outputs[3] [24]), 
         .C(n23465), .D(n2022[17]), .Z(n66354)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_275.init = 16'hfefa;
    LUT4 i1_4_lut_adj_276 (.A(\hidden_outputs[3] [23]), .B(n22568), .C(float_alu_c[23]), 
         .D(n70785), .Z(n22694)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_276.init = 16'hc088;
    LUT4 i2_4_lut_adj_277 (.A(n10_adj_191), .B(n22694), .C(\hidden_outputs[3] [23]), 
         .D(n2022[17]), .Z(n62938)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_277.init = 16'hfeee;
    LUT4 i1_4_lut_adj_278 (.A(\hidden_outputs[3] [22]), .B(n22568), .C(float_alu_c[22]), 
         .D(n70785), .Z(n23459)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_278.init = 16'hc088;
    LUT4 i1_4_lut_adj_279 (.A(n10_adj_192), .B(\hidden_outputs[3] [22]), 
         .C(n23459), .D(n2022[17]), .Z(n66358)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_279.init = 16'hfefa;
    LUT4 i1_4_lut_adj_280 (.A(\hidden_outputs[3] [21]), .B(n22568), .C(float_alu_c[21]), 
         .D(n70785), .Z(n22697)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_280.init = 16'hc088;
    LUT4 i12598_2_lut_4_lut_3_lut (.A(n2022[38]), .B(n70822), .C(n2022[31]), 
         .Z(n24288)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i12598_2_lut_4_lut_3_lut.init = 16'h4040;
    LUT4 i2_4_lut_adj_281 (.A(n10_adj_193), .B(n22697), .C(\hidden_outputs[3] [21]), 
         .D(n2022[17]), .Z(n62940)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_281.init = 16'hfeee;
    LUT4 i1_4_lut_adj_282 (.A(\hidden_outputs[3] [20]), .B(n22568), .C(float_alu_c[20]), 
         .D(n70785), .Z(n23417)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_282.init = 16'hc088;
    LUT4 i1_4_lut_adj_283 (.A(n10_adj_194), .B(\hidden_outputs[3] [20]), 
         .C(n23417), .D(n2022[17]), .Z(n66496)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_283.init = 16'hfefa;
    LUT4 i1_4_lut_adj_284 (.A(\hidden_outputs[3] [19]), .B(n22568), .C(float_alu_c[19]), 
         .D(n70785), .Z(n22700)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_284.init = 16'hc088;
    PFUMX i54520 (.BLUT(n67429), .ALUT(n67430), .C0(h[1]), .Z(n67431));
    LUT4 i1_4_lut_adj_285 (.A(n10_adj_195), .B(n22700), .C(\hidden_outputs[3] [19]), 
         .D(n2022[17]), .Z(n66482)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_285.init = 16'hfeee;
    PFUMX i54523 (.BLUT(n67432), .ALUT(n67433), .C0(h[1]), .Z(n67434));
    LUT4 i1_4_lut_adj_286 (.A(\hidden_outputs[3] [18]), .B(n22568), .C(float_alu_c[18]), 
         .D(n70785), .Z(n23405)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_286.init = 16'hc088;
    LUT4 i1_4_lut_adj_287 (.A(n10_adj_196), .B(\hidden_outputs[3] [18]), 
         .C(n23405), .D(n2022[17]), .Z(n66372)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_287.init = 16'hfefa;
    PFUMX i54526 (.BLUT(n67435), .ALUT(n67436), .C0(h[1]), .Z(n67437));
    LUT4 i1_4_lut_adj_288 (.A(\hidden_outputs[3] [17]), .B(n22568), .C(float_alu_c[17]), 
         .D(n70785), .Z(n22703)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_288.init = 16'hc088;
    PFUMX i54529 (.BLUT(n67438), .ALUT(n67439), .C0(h[1]), .Z(n67440));
    LUT4 i2_4_lut_adj_289 (.A(n10_adj_199), .B(n22703), .C(\hidden_outputs[3] [17]), 
         .D(n2022[17]), .Z(n62942)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_289.init = 16'hfeee;
    LUT4 i1_4_lut_adj_290 (.A(\hidden_outputs[3] [16]), .B(n22568), .C(float_alu_c[16]), 
         .D(n70785), .Z(n23390)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_290.init = 16'hc088;
    PFUMX i54532 (.BLUT(n67441), .ALUT(n67442), .C0(h[1]), .Z(n67443));
    LUT4 i2_4_lut_adj_291 (.A(n23390), .B(n10_adj_205), .C(\hidden_outputs[3] [16]), 
         .D(n2022[17]), .Z(n63199)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_291.init = 16'hfeee;
    PFUMX i54535 (.BLUT(n67444), .ALUT(n67445), .C0(h[1]), .Z(n67446));
    PFUMX i54538 (.BLUT(n67447), .ALUT(n67448), .C0(h[1]), .Z(n67449));
    LUT4 i1_4_lut_adj_292 (.A(\hidden_outputs[3] [15]), .B(n22568), .C(float_alu_c[15]), 
         .D(n70785), .Z(n22706)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_292.init = 16'hc088;
    LUT4 i1_4_lut_adj_293 (.A(n10_adj_207), .B(n22706), .C(\hidden_outputs[3] [15]), 
         .D(n2022[17]), .Z(n66480)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_293.init = 16'hfeee;
    LUT4 i1_4_lut_adj_294 (.A(\hidden_outputs[3] [14]), .B(n22568), .C(float_alu_c[14]), 
         .D(n70785), .Z(n23315)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_294.init = 16'hc088;
    PFUMX i54541 (.BLUT(n67450), .ALUT(n67451), .C0(n[1]), .Z(n67452));
    LUT4 i1_4_lut_adj_295 (.A(n10_adj_222), .B(\hidden_outputs[3] [14]), 
         .C(n23315), .D(n2022[17]), .Z(n66554)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_295.init = 16'hfefa;
    PFUMX i54544 (.BLUT(n67453), .ALUT(n67454), .C0(n[1]), .Z(n67455));
    PFUMX i54547 (.BLUT(n67456), .ALUT(n67457), .C0(n[1]), .Z(n67458));
    PFUMX i54550 (.BLUT(n67459), .ALUT(n67460), .C0(n[1]), .Z(n67461));
    PFUMX i54553 (.BLUT(n67462), .ALUT(n67463), .C0(n[1]), .Z(n67464));
    LUT4 i1_4_lut_adj_296 (.A(\hidden_outputs[3] [13]), .B(n22568), .C(float_alu_c[13]), 
         .D(n70785), .Z(n23312)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_296.init = 16'hc088;
    LUT4 i2_4_lut_adj_297 (.A(n23312), .B(n10_adj_224), .C(\hidden_outputs[3] [13]), 
         .D(n2022[17]), .Z(n63173)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_297.init = 16'hfeee;
    FD1P3DX done_438 (.D(n3756), .SP(n77), .CK(clock), .CD(SDA_c), .Q(mlp_done));
    defparam done_438.GSR = "DISABLED";
    FD1P3BX state_FSM__i1 (.D(n73801), .SP(n64), .CK(clock), .PD(SDA_c), 
            .Q(n2086));
    defparam state_FSM__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_298 (.A(\hidden_outputs[3] [12]), .B(n22568), .C(float_alu_c[12]), 
         .D(n70785), .Z(n22712)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_298.init = 16'hc088;
    LUT4 i2_4_lut_adj_299 (.A(n10_adj_225), .B(n22712), .C(\hidden_outputs[3] [12]), 
         .D(n2022[17]), .Z(n62944)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_299.init = 16'hfeee;
    LUT4 i1_4_lut_adj_300 (.A(\hidden_outputs[3] [11]), .B(n22568), .C(float_alu_c[11]), 
         .D(n70785), .Z(n23309)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_300.init = 16'hc088;
    LUT4 i1_4_lut_adj_301 (.A(n10_adj_226), .B(\hidden_outputs[3] [11]), 
         .C(n23309), .D(n2022[17]), .Z(n66392)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_301.init = 16'hfefa;
    LUT4 i1_4_lut_adj_302 (.A(\hidden_outputs[3] [10]), .B(n22568), .C(float_alu_c[10]), 
         .D(n70785), .Z(n22715)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_302.init = 16'hc088;
    LUT4 i1_4_lut_adj_303 (.A(n10_adj_227), .B(n22715), .C(\hidden_outputs[3] [10]), 
         .D(n2022[17]), .Z(n66478)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_303.init = 16'hfeee;
    LUT4 i1_4_lut_adj_304 (.A(\hidden_outputs[3] [9]), .B(n22568), .C(float_alu_c[9]), 
         .D(n70785), .Z(n23306)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_304.init = 16'hc088;
    LUT4 i1_4_lut_adj_305 (.A(n10_adj_228), .B(\hidden_outputs[3] [9]), 
         .C(n23306), .D(n2022[17]), .Z(n66552)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_305.init = 16'hfefa;
    LUT4 i1_4_lut_adj_306 (.A(\hidden_outputs[3] [8]), .B(n22568), .C(float_alu_c[8]), 
         .D(n70785), .Z(n23303)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_306.init = 16'hc088;
    LUT4 i1_4_lut_adj_307 (.A(n10_adj_229), .B(\hidden_outputs[3] [8]), 
         .C(n23303), .D(n2022[17]), .Z(n66394)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_307.init = 16'hfefa;
    LUT4 i1_4_lut_adj_308 (.A(\hidden_outputs[3] [7]), .B(n22568), .C(float_alu_c[7]), 
         .D(n70785), .Z(n22718)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_308.init = 16'hc088;
    LUT4 i2_4_lut_adj_309 (.A(n10_adj_230), .B(n22718), .C(\hidden_outputs[3] [7]), 
         .D(n2022[17]), .Z(n62946)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_309.init = 16'hfeee;
    LUT4 i1_4_lut_adj_310 (.A(\hidden_outputs[3] [6]), .B(n22568), .C(float_alu_c[6]), 
         .D(n70785), .Z(n23300)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_310.init = 16'hc088;
    LUT4 i2_4_lut_adj_311 (.A(n23300), .B(n10_adj_231), .C(\hidden_outputs[3] [6]), 
         .D(n2022[17]), .Z(n63168)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_311.init = 16'hfeee;
    LUT4 i1_4_lut_adj_312 (.A(\hidden_outputs[3] [5]), .B(n22568), .C(float_alu_c[5]), 
         .D(n70785), .Z(n22721)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_312.init = 16'hc088;
    LUT4 i1_4_lut_adj_313 (.A(n10_adj_232), .B(n22721), .C(\hidden_outputs[3] [5]), 
         .D(n2022[17]), .Z(n66476)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_313.init = 16'hfeee;
    LUT4 i1_4_lut_adj_314 (.A(\hidden_outputs[3] [4]), .B(n22568), .C(float_alu_c[4]), 
         .D(n70785), .Z(n22724)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_314.init = 16'hc088;
    LUT4 i2_4_lut_adj_315 (.A(n10_adj_233), .B(n22724), .C(\hidden_outputs[3] [4]), 
         .D(n2022[17]), .Z(n62948)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_315.init = 16'hfeee;
    LUT4 i1_4_lut_adj_316 (.A(\hidden_outputs[3] [3]), .B(n22568), .C(float_alu_c[3]), 
         .D(n70785), .Z(n22727)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_316.init = 16'hc088;
    LUT4 i2_4_lut_adj_317 (.A(n10_adj_234), .B(n22727), .C(\hidden_outputs[3] [3]), 
         .D(n2022[17]), .Z(n62949)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_317.init = 16'hfeee;
    LUT4 i1_4_lut_adj_318 (.A(\hidden_outputs[3] [2]), .B(n22568), .C(float_alu_c[2]), 
         .D(n70785), .Z(n23291)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_318.init = 16'hc088;
    LUT4 i1_4_lut_adj_319 (.A(n10_adj_235), .B(\hidden_outputs[3] [2]), 
         .C(n23291), .D(n2022[17]), .Z(n66486)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_319.init = 16'hfefa;
    LUT4 i1_4_lut_adj_320 (.A(\hidden_outputs[3] [1]), .B(n22568), .C(float_alu_c[1]), 
         .D(n70785), .Z(n22730)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_320.init = 16'hc088;
    LUT4 i1_4_lut_adj_321 (.A(n10_adj_236), .B(n22730), .C(\hidden_outputs[3] [1]), 
         .D(n2022[17]), .Z(n66472)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_321.init = 16'hfeee;
    LUT4 i54489_3_lut (.A(\hidden_outputs[2] [15]), .B(\hidden_outputs[3] [15]), 
         .C(h[0]), .Z(n67400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54489_3_lut.init = 16'hcaca;
    LUT4 i54488_3_lut (.A(\hidden_outputs[0] [15]), .B(\hidden_outputs[1] [15]), 
         .C(h[0]), .Z(n67399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54488_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_322 (.A(\state[0] ), .B(n3946), .C(n3944), .D(weight_done), 
         .Z(n22106)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_322.init = 16'hfaee;
    LUT4 i34469_3_lut (.A(n3944), .B(n3946), .C(weight_done), .Z(n3961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i34469_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_323 (.A(\hidden_outputs[2] [31]), .B(n22568), .C(float_alu_c[31]), 
         .D(n70787), .Z(n22637)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_323.init = 16'hc088;
    LUT4 i1_4_lut_adj_324 (.A(n10_adj_182), .B(n22637), .C(n1584), .D(n2022[17]), 
         .Z(n66512)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_324.init = 16'hfeee;
    LUT4 i1_4_lut_adj_325 (.A(\hidden_outputs[2] [30]), .B(n22568), .C(float_alu_c[30]), 
         .D(n70787), .Z(n23270)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_325.init = 16'hc088;
    LUT4 i2_4_lut_adj_326 (.A(n23270), .B(n10_adj_183), .C(\hidden_outputs[2] [30]), 
         .D(n2022[17]), .Z(n63080)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_326.init = 16'hfeee;
    LUT4 i1_4_lut_adj_327 (.A(\hidden_outputs[2] [29]), .B(n22568), .C(float_alu_c[29]), 
         .D(n70787), .Z(n22640)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_327.init = 16'hc088;
    LUT4 i2_4_lut_adj_328 (.A(n10_adj_185), .B(n22640), .C(\hidden_outputs[2] [29]), 
         .D(n2022[17]), .Z(n62914)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_328.init = 16'hfeee;
    LUT4 i1_4_lut_adj_329 (.A(\hidden_outputs[2] [28]), .B(n22568), .C(float_alu_c[28]), 
         .D(n70787), .Z(n23267)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_329.init = 16'hc088;
    LUT4 i1_4_lut_adj_330 (.A(n10_adj_186), .B(\hidden_outputs[2] [28]), 
         .C(n23267), .D(n2022[17]), .Z(n66266)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_330.init = 16'hfefa;
    LUT4 i1_4_lut_adj_331 (.A(\hidden_outputs[2] [27]), .B(n22568), .C(float_alu_c[27]), 
         .D(n70787), .Z(n23264)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_331.init = 16'hc088;
    LUT4 i1_4_lut_adj_332 (.A(n10_adj_187), .B(\hidden_outputs[2] [27]), 
         .C(n23264), .D(n2022[17]), .Z(n66288)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_332.init = 16'hfefa;
    LUT4 i1_4_lut_adj_333 (.A(\hidden_outputs[2] [26]), .B(n22568), .C(float_alu_c[26]), 
         .D(n70787), .Z(n22643)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_333.init = 16'hc088;
    LUT4 i1_4_lut_adj_334 (.A(n10_adj_188), .B(n22643), .C(\hidden_outputs[2] [26]), 
         .D(n2022[17]), .Z(n66510)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_334.init = 16'hfeee;
    LUT4 i1_4_lut_adj_335 (.A(\hidden_outputs[2] [25]), .B(n22568), .C(float_alu_c[25]), 
         .D(n70787), .Z(n23258)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_335.init = 16'hc088;
    LUT4 i2_4_lut_adj_336 (.A(n23258), .B(n10_adj_189), .C(\hidden_outputs[2] [25]), 
         .D(n2022[17]), .Z(n63085)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_336.init = 16'hfeee;
    LUT4 i1_4_lut_adj_337 (.A(\hidden_outputs[2] [24]), .B(n22568), .C(float_alu_c[24]), 
         .D(n70787), .Z(n22646)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_337.init = 16'hc088;
    LUT4 i2_4_lut_adj_338 (.A(n10_adj_190), .B(n22646), .C(\hidden_outputs[2] [24]), 
         .D(n2022[17]), .Z(n62916)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_338.init = 16'hfeee;
    LUT4 i1_4_lut_adj_339 (.A(\hidden_outputs[2] [23]), .B(n22568), .C(float_alu_c[23]), 
         .D(n70787), .Z(n23255)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_339.init = 16'hc088;
    LUT4 i1_4_lut_adj_340 (.A(n10_adj_191), .B(\hidden_outputs[2] [23]), 
         .C(n23255), .D(n2022[17]), .Z(n66294)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_340.init = 16'hfefa;
    LUT4 i1_4_lut_adj_341 (.A(\hidden_outputs[2] [22]), .B(n22568), .C(float_alu_c[22]), 
         .D(n70787), .Z(n22649)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_341.init = 16'hc088;
    LUT4 i1_4_lut_adj_342 (.A(n10_adj_192), .B(n22649), .C(\hidden_outputs[2] [22]), 
         .D(n2022[17]), .Z(n66508)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_342.init = 16'hfeee;
    LUT4 i1_4_lut_adj_343 (.A(\hidden_outputs[2] [21]), .B(n22568), .C(float_alu_c[21]), 
         .D(n70787), .Z(n23252)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_343.init = 16'hc088;
    PFUMX i54556 (.BLUT(n67465), .ALUT(n67466), .C0(n[1]), .Z(n67467));
    LUT4 i2_4_lut_adj_344 (.A(n23252), .B(n10_adj_193), .C(\hidden_outputs[2] [21]), 
         .D(n2022[17]), .Z(n63078)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_344.init = 16'hfeee;
    LUT4 i1_4_lut_adj_345 (.A(\hidden_outputs[2] [20]), .B(n22568), .C(float_alu_c[20]), 
         .D(n70787), .Z(n22652)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_345.init = 16'hc088;
    LUT4 i1_4_lut_adj_346 (.A(n10_adj_194), .B(n22652), .C(\hidden_outputs[2] [20]), 
         .D(n2022[17]), .Z(n66406)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_346.init = 16'hfeee;
    PFUMX i54559 (.BLUT(n67468), .ALUT(n67469), .C0(n[1]), .Z(n67470));
    LUT4 i1_4_lut_adj_347 (.A(\hidden_outputs[2] [19]), .B(n22568), .C(float_alu_c[19]), 
         .D(n70787), .Z(n23246)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_347.init = 16'hc088;
    LUT4 i1_4_lut_adj_348 (.A(n10_adj_195), .B(\hidden_outputs[2] [19]), 
         .C(n23246), .D(n2022[17]), .Z(n66290)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_348.init = 16'hfefa;
    LUT4 i1_4_lut_adj_349 (.A(\hidden_outputs[2] [18]), .B(n22568), .C(float_alu_c[18]), 
         .D(n70787), .Z(n22655)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_349.init = 16'hc088;
    LUT4 i2_4_lut_adj_350 (.A(n10_adj_196), .B(n22655), .C(\hidden_outputs[2] [18]), 
         .D(n2022[17]), .Z(n62920)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_350.init = 16'hfeee;
    LUT4 i1_4_lut_adj_351 (.A(\hidden_outputs[2] [17]), .B(n22568), .C(float_alu_c[17]), 
         .D(n70787), .Z(n23243)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_351.init = 16'hc088;
    PFUMX i54562 (.BLUT(n67471), .ALUT(n67472), .C0(n[1]), .Z(n67473));
    LUT4 i2_4_lut_adj_352 (.A(n23243), .B(n10_adj_199), .C(\hidden_outputs[2] [17]), 
         .D(n2022[17]), .Z(n63083)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_352.init = 16'hfeee;
    LUT4 i1_4_lut_adj_353 (.A(\hidden_outputs[2] [16]), .B(n22568), .C(float_alu_c[16]), 
         .D(n70787), .Z(n22658)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_353.init = 16'hc088;
    PFUMX i54565 (.BLUT(n67474), .ALUT(n67475), .C0(n[1]), .Z(n67476));
    LUT4 i1_4_lut_adj_354 (.A(n10_adj_205), .B(n22658), .C(\hidden_outputs[2] [16]), 
         .D(n2022[17]), .Z(n66506)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_354.init = 16'hfeee;
    LUT4 i1_4_lut_adj_355 (.A(\hidden_outputs[2] [15]), .B(n22568), .C(float_alu_c[15]), 
         .D(n70787), .Z(n23372)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_355.init = 16'hc088;
    FD1P3IX numL_4656__i0 (.D(n134_adj_407[0]), .SP(n70817), .CD(n24021), 
            .CK(clock), .Q(numL[0]));
    defparam numL_4656__i0.GSR = "DISABLED";
    PFUMX i54568 (.BLUT(n67477), .ALUT(n67478), .C0(n[1]), .Z(n67479));
    LUT4 i2_4_lut_adj_356 (.A(n23372), .B(n10_adj_207), .C(\hidden_outputs[2] [15]), 
         .D(n2022[17]), .Z(n63192)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_356.init = 16'hfeee;
    PFUMX i54571 (.BLUT(n67480), .ALUT(n67481), .C0(n[1]), .Z(n67482));
    LUT4 i1_4_lut_adj_357 (.A(\hidden_outputs[2] [14]), .B(n22568), .C(float_alu_c[14]), 
         .D(n70787), .Z(n23231)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_357.init = 16'hc088;
    LUT4 i1_4_lut_adj_358 (.A(n10_adj_222), .B(\hidden_outputs[2] [14]), 
         .C(n23231), .D(n2022[17]), .Z(n66274)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_358.init = 16'hfefa;
    LUT4 i1_4_lut_adj_359 (.A(\hidden_outputs[2] [13]), .B(n22568), .C(float_alu_c[13]), 
         .D(n70787), .Z(n22661)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_359.init = 16'hc088;
    LUT4 i2_4_lut_adj_360 (.A(n10_adj_224), .B(n22661), .C(\hidden_outputs[2] [13]), 
         .D(n2022[17]), .Z(n62922)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_360.init = 16'hfeee;
    LUT4 i1_4_lut_adj_361 (.A(\hidden_outputs[2] [12]), .B(n22568), .C(float_alu_c[12]), 
         .D(n70787), .Z(n23228)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_361.init = 16'hc088;
    LUT4 i1_4_lut_adj_362 (.A(n10_adj_225), .B(\hidden_outputs[2] [12]), 
         .C(n23228), .D(n2022[17]), .Z(n66272)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_362.init = 16'hfefa;
    LUT4 i1_4_lut_adj_363 (.A(\hidden_outputs[2] [11]), .B(n22568), .C(float_alu_c[11]), 
         .D(n70787), .Z(n22664)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_363.init = 16'hc088;
    LUT4 i1_4_lut_adj_364 (.A(n10_adj_226), .B(n22664), .C(\hidden_outputs[2] [11]), 
         .D(n2022[17]), .Z(n66504)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_364.init = 16'hfeee;
    LUT4 i1_4_lut_adj_365 (.A(\hidden_outputs[2] [10]), .B(n22568), .C(float_alu_c[10]), 
         .D(n70787), .Z(n23225)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_365.init = 16'hc088;
    LUT4 i2_4_lut_adj_366 (.A(n23225), .B(n10_adj_227), .C(\hidden_outputs[2] [10]), 
         .D(n2022[17]), .Z(n63091)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_366.init = 16'hfeee;
    LUT4 i1_4_lut_adj_367 (.A(\hidden_outputs[2] [9]), .B(n22568), .C(float_alu_c[9]), 
         .D(n70787), .Z(n23222)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_367.init = 16'hc088;
    LUT4 i1_4_lut_adj_368 (.A(n10_adj_228), .B(\hidden_outputs[2] [9]), 
         .C(n23222), .D(n2022[17]), .Z(n66304)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_368.init = 16'hfefa;
    LUT4 i1_4_lut_adj_369 (.A(\hidden_outputs[2] [8]), .B(n22568), .C(float_alu_c[8]), 
         .D(n70787), .Z(n22667)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_369.init = 16'hc088;
    LUT4 i1_4_lut_adj_370 (.A(n10_adj_229), .B(n22667), .C(\hidden_outputs[2] [8]), 
         .D(n2022[17]), .Z(n66502)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_370.init = 16'hfeee;
    LUT4 i1_4_lut_adj_371 (.A(\hidden_outputs[2] [7]), .B(n22568), .C(float_alu_c[7]), 
         .D(n70787), .Z(n22670)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_371.init = 16'hc088;
    LUT4 i2_4_lut_adj_372 (.A(n10_adj_230), .B(n22670), .C(\hidden_outputs[2] [7]), 
         .D(n2022[17]), .Z(n62925)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_372.init = 16'hfeee;
    LUT4 i1_4_lut_adj_373 (.A(\hidden_outputs[2] [6]), .B(n22568), .C(float_alu_c[6]), 
         .D(n70787), .Z(n23210)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_373.init = 16'hc088;
    LUT4 i2_4_lut_adj_374 (.A(n23210), .B(n10_adj_231), .C(\hidden_outputs[2] [6]), 
         .D(n2022[17]), .Z(n63094)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_374.init = 16'hfeee;
    LUT4 i1_4_lut_adj_375 (.A(\hidden_outputs[2] [5]), .B(n22568), .C(float_alu_c[5]), 
         .D(n70787), .Z(n22673)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_375.init = 16'hc088;
    LUT4 i1_4_lut_adj_376 (.A(n10_adj_232), .B(n22673), .C(\hidden_outputs[2] [5]), 
         .D(n2022[17]), .Z(n66500)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_376.init = 16'hfeee;
    LUT4 i1_4_lut_adj_377 (.A(\hidden_outputs[2] [4]), .B(n22568), .C(float_alu_c[4]), 
         .D(n70787), .Z(n23201)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_377.init = 16'hc088;
    LUT4 i2_4_lut_adj_378 (.A(n23201), .B(n10_adj_233), .C(\hidden_outputs[2] [4]), 
         .D(n2022[17]), .Z(n63093)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_378.init = 16'hfeee;
    LUT4 i1_4_lut_adj_379 (.A(\hidden_outputs[2] [3]), .B(n22568), .C(float_alu_c[3]), 
         .D(n70787), .Z(n22676)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_379.init = 16'hc088;
    LUT4 i1_4_lut_adj_380 (.A(n10_adj_234), .B(n22676), .C(\hidden_outputs[2] [3]), 
         .D(n2022[17]), .Z(n66492)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_380.init = 16'hfeee;
    LUT4 i1_4_lut_adj_381 (.A(\hidden_outputs[2] [2]), .B(n22568), .C(float_alu_c[2]), 
         .D(n70787), .Z(n22679)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_381.init = 16'hc088;
    FD1P3IX h_4657__i0 (.D(n134[0]), .SP(n23680), .CD(n24020), .CK(clock), 
            .Q(h[0]));
    defparam h_4657__i0.GSR = "DISABLED";
    FD1P3IX n_4659__i29 (.D(n134_adj_403[29]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[29]));
    defparam n_4659__i29.GSR = "DISABLED";
    FD1P3IX n_4659__i0 (.D(n134_adj_403[0]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[0]));
    defparam n_4659__i0.GSR = "DISABLED";
    LUT4 i2_4_lut_adj_382 (.A(n10_adj_235), .B(n22679), .C(\hidden_outputs[2] [2]), 
         .D(n2022[17]), .Z(n62932)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_382.init = 16'hfeee;
    LUT4 i1_4_lut_adj_383 (.A(\hidden_outputs[2] [1]), .B(n22568), .C(float_alu_c[1]), 
         .D(n70787), .Z(n23195)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_383.init = 16'hc088;
    CCU2D equal_232_32 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n60990), 
          .S0(n3922));
    defparam equal_232_32.INIT0 = 16'hFFFF;
    defparam equal_232_32.INIT1 = 16'h0000;
    defparam equal_232_32.INJECT1_0 = "NO";
    defparam equal_232_32.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_384 (.A(n10_adj_236), .B(\hidden_outputs[2] [1]), 
         .C(n23195), .D(n2022[17]), .Z(n66296)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_384.init = 16'hfefa;
    LUT4 i1_4_lut_adj_385 (.A(\hidden_outputs[1] [31]), .B(n22568), .C(float_alu_c[31]), 
         .D(n70789), .Z(n22598)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_385.init = 16'hc088;
    LUT4 i1_4_lut_adj_386 (.A(n10_adj_182), .B(n22598), .C(n1585), .D(n2022[17]), 
         .Z(n66324)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_386.init = 16'hfeee;
    LUT4 i1_4_lut_adj_387 (.A(\hidden_outputs[1] [30]), .B(n22568), .C(float_alu_c[30]), 
         .D(n70789), .Z(n22874)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_387.init = 16'hc088;
    LUT4 i1_4_lut_adj_388 (.A(n10_adj_183), .B(n22874), .C(\hidden_outputs[1] [30]), 
         .D(n2022[17]), .Z(n66430)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_388.init = 16'hfeee;
    LUT4 i1_4_lut_adj_389 (.A(\hidden_outputs[1] [29]), .B(n22568), .C(float_alu_c[29]), 
         .D(n70789), .Z(n22601)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_389.init = 16'hc088;
    PFUMX i54574 (.BLUT(n67483), .ALUT(n67484), .C0(n[1]), .Z(n67485));
    PFUMX i54577 (.BLUT(n67486), .ALUT(n67487), .C0(n[1]), .Z(n67488));
    PFUMX i54580 (.BLUT(n67489), .ALUT(n67490), .C0(n[1]), .Z(n67491));
    PFUMX i54583 (.BLUT(n67492), .ALUT(n67493), .C0(n[1]), .Z(n67494));
    LUT4 i2_4_lut_adj_390 (.A(n10_adj_185), .B(n22601), .C(\hidden_outputs[1] [29]), 
         .D(n2022[17]), .Z(n62899)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_390.init = 16'hfeee;
    PFUMX i54586 (.BLUT(n67495), .ALUT(n67496), .C0(n[1]), .Z(n67497));
    PFUMX i54589 (.BLUT(n67498), .ALUT(n67499), .C0(n[1]), .Z(n67500));
    LUT4 i1_4_lut_adj_391 (.A(\hidden_outputs[1] [28]), .B(n22568), .C(float_alu_c[28]), 
         .D(n70789), .Z(n22841)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_391.init = 16'hc088;
    PFUMX i54592 (.BLUT(n67501), .ALUT(n67502), .C0(n[1]), .Z(n67503));
    PFUMX i54595 (.BLUT(n67504), .ALUT(n67505), .C0(n[1]), .Z(n67506));
    PFUMX i54598 (.BLUT(n67507), .ALUT(n67508), .C0(n[1]), .Z(n67509));
    LUT4 i1_4_lut_adj_392 (.A(n10_adj_186), .B(\hidden_outputs[1] [28]), 
         .C(n22841), .D(n2022[17]), .Z(n66332)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_392.init = 16'hfefa;
    LUT4 i1_4_lut_adj_393 (.A(\hidden_outputs[1] [27]), .B(n22568), .C(float_alu_c[27]), 
         .D(n70789), .Z(n22898)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_393.init = 16'hc088;
    FD1P3IX n_4659__i28 (.D(n134_adj_403[28]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[28]));
    defparam n_4659__i28.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_394 (.A(n10_adj_187), .B(n22898), .C(\hidden_outputs[1] [27]), 
         .D(n2022[17]), .Z(n66418)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_394.init = 16'hfeee;
    LUT4 i1_4_lut_adj_395 (.A(\hidden_outputs[1] [26]), .B(n22568), .C(float_alu_c[26]), 
         .D(n70789), .Z(n23387)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_395.init = 16'hc088;
    LUT4 i1_4_lut_adj_396 (.A(n10_adj_188), .B(\hidden_outputs[1] [26]), 
         .C(n23387), .D(n2022[17]), .Z(n66378)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_396.init = 16'hfefa;
    LUT4 i1_4_lut_adj_397 (.A(\hidden_outputs[1] [25]), .B(n22568), .C(float_alu_c[25]), 
         .D(n70789), .Z(n22901)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_397.init = 16'hc088;
    PFUMX i54601 (.BLUT(n67510), .ALUT(n67511), .C0(n[1]), .Z(n67512));
    LUT4 i2_4_lut_adj_398 (.A(n10_adj_189), .B(n22901), .C(\hidden_outputs[1] [25]), 
         .D(n2022[17]), .Z(n63004)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_398.init = 16'hfeee;
    LUT4 i1_4_lut_adj_399 (.A(\hidden_outputs[1] [24]), .B(n22568), .C(float_alu_c[24]), 
         .D(n70789), .Z(n23384)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_399.init = 16'hc088;
    LUT4 i2_4_lut_adj_400 (.A(n23384), .B(n10_adj_190), .C(\hidden_outputs[1] [24]), 
         .D(n2022[17]), .Z(n63197)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_400.init = 16'hfeee;
    LUT4 i1_4_lut_adj_401 (.A(\hidden_outputs[1] [23]), .B(n22568), .C(float_alu_c[23]), 
         .D(n70789), .Z(n22904)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_401.init = 16'hc088;
    LUT4 i1_4_lut_adj_402 (.A(n10_adj_191), .B(n22904), .C(\hidden_outputs[1] [23]), 
         .D(n2022[17]), .Z(n66416)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_402.init = 16'hfeee;
    LUT4 i1_4_lut_adj_403 (.A(\hidden_outputs[1] [22]), .B(n22568), .C(float_alu_c[22]), 
         .D(n70789), .Z(n23381)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_403.init = 16'hc088;
    FD1P3IX n_4659__i27 (.D(n134_adj_403[27]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[27]));
    defparam n_4659__i27.GSR = "DISABLED";
    FD1P3IX o_4661__i0 (.D(n134_adj_404[0]), .SP(n73800), .CD(n24257), 
            .CK(clock), .Q(o[0]));
    defparam o_4661__i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_404 (.A(n10_adj_192), .B(\hidden_outputs[1] [22]), 
         .C(n23381), .D(n2022[17]), .Z(n66380)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_404.init = 16'hfefa;
    LUT4 i1_4_lut_adj_405 (.A(\hidden_outputs[1] [21]), .B(n22568), .C(float_alu_c[21]), 
         .D(n70789), .Z(n22907)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_405.init = 16'hc088;
    LUT4 i1_4_lut_adj_406 (.A(n10_adj_193), .B(n22907), .C(\hidden_outputs[1] [21]), 
         .D(n2022[17]), .Z(n66414)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_406.init = 16'hfeee;
    LUT4 i1_4_lut_adj_407 (.A(\hidden_outputs[1] [20]), .B(n22568), .C(float_alu_c[20]), 
         .D(n70789), .Z(n23378)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_407.init = 16'hc088;
    LUT4 i2_4_lut_adj_408 (.A(n23378), .B(n10_adj_194), .C(\hidden_outputs[1] [20]), 
         .D(n2022[17]), .Z(n63194)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_408.init = 16'hfeee;
    LUT4 i1_4_lut_adj_409 (.A(\hidden_outputs[1] [19]), .B(n22568), .C(float_alu_c[19]), 
         .D(n70789), .Z(n23375)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_409.init = 16'hc088;
    LUT4 i1_4_lut_adj_410 (.A(n10_adj_195), .B(\hidden_outputs[1] [19]), 
         .C(n23375), .D(n2022[17]), .Z(n66382)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_410.init = 16'hfefa;
    LUT4 i1_4_lut_adj_411 (.A(\hidden_outputs[1] [18]), .B(n22568), .C(float_alu_c[18]), 
         .D(n70789), .Z(n23420)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_411.init = 16'hc088;
    LUT4 i1_4_lut_adj_412 (.A(n10_adj_196), .B(\hidden_outputs[1] [18]), 
         .C(n23420), .D(n2022[17]), .Z(n66370)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_412.init = 16'hfefa;
    LUT4 i1_4_lut_adj_413 (.A(\hidden_outputs[1] [17]), .B(n22568), .C(float_alu_c[17]), 
         .D(n70789), .Z(n22826)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_413.init = 16'hc088;
    LUT4 i1_4_lut_adj_414 (.A(n10_adj_199), .B(\hidden_outputs[1] [17]), 
         .C(n22826), .D(n2022[17]), .Z(n66308)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_414.init = 16'hfefa;
    LUT4 i1_4_lut_adj_415 (.A(\hidden_outputs[1] [16]), .B(n22568), .C(float_alu_c[16]), 
         .D(n70789), .Z(n22910)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_415.init = 16'hc088;
    LUT4 i1_4_lut_adj_416 (.A(n10_adj_205), .B(n22910), .C(\hidden_outputs[1] [16]), 
         .D(n2022[17]), .Z(n66410)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_416.init = 16'hfeee;
    FD1P3IX n_4659__i26 (.D(n134_adj_403[26]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[26]));
    defparam n_4659__i26.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_417 (.A(\hidden_outputs[1] [15]), .B(n22568), .C(float_alu_c[15]), 
         .D(n70789), .Z(n22613)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_417.init = 16'hc088;
    PFUMX i54604 (.BLUT(n67513), .ALUT(n67514), .C0(n[1]), .Z(n67515));
    FD1P3IX n_4659__i25 (.D(n134_adj_403[25]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[25]));
    defparam n_4659__i25.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_418 (.A(n10_adj_207), .B(n22613), .C(\hidden_outputs[1] [15]), 
         .D(n2022[17]), .Z(n66520)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_418.init = 16'hfeee;
    FD1P3IX n_4659__i24 (.D(n134_adj_403[24]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[24]));
    defparam n_4659__i24.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_419 (.A(\hidden_outputs[1] [14]), .B(n22568), .C(float_alu_c[14]), 
         .D(n70789), .Z(n22616)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_419.init = 16'hc088;
    FD1P3IX n_4659__i23 (.D(n134_adj_403[23]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[23]));
    defparam n_4659__i23.GSR = "DISABLED";
    LUT4 i2_4_lut_adj_420 (.A(n10_adj_222), .B(n22616), .C(\hidden_outputs[1] [14]), 
         .D(n2022[17]), .Z(n62905)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_420.init = 16'hfeee;
    FD1P3IX n_4659__i22 (.D(n134_adj_403[22]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[22]));
    defparam n_4659__i22.GSR = "DISABLED";
    PFUMX i54607 (.BLUT(n67516), .ALUT(n67517), .C0(n[1]), .Z(n67518));
    PFUMX i54610 (.BLUT(n67519), .ALUT(n67520), .C0(n[1]), .Z(n67521));
    LUT4 i1_4_lut_adj_421 (.A(\hidden_outputs[1] [13]), .B(n22568), .C(float_alu_c[13]), 
         .D(n70789), .Z(n22709)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_421.init = 16'hc088;
    LUT4 i1_4_lut_adj_422 (.A(n10_adj_224), .B(\hidden_outputs[1] [13]), 
         .C(n22709), .D(n2022[17]), .Z(n66562)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_422.init = 16'hfefa;
    LUT4 i1_4_lut_adj_423 (.A(\hidden_outputs[1] [12]), .B(n22568), .C(float_alu_c[12]), 
         .D(n70789), .Z(n22619)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_423.init = 16'hc088;
    LUT4 i1_4_lut_adj_424 (.A(n10_adj_225), .B(n22619), .C(\hidden_outputs[1] [12]), 
         .D(n2022[17]), .Z(n66518)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_424.init = 16'hfeee;
    LUT4 i1_4_lut_adj_425 (.A(\hidden_outputs[1] [11]), .B(n22568), .C(float_alu_c[11]), 
         .D(n70789), .Z(n22583)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_425.init = 16'hc088;
    LUT4 i1_4_lut_adj_426 (.A(n10_adj_226), .B(\hidden_outputs[1] [11]), 
         .C(n22583), .D(n2022[17]), .Z(n66314)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_426.init = 16'hfefa;
    LUT4 i1_4_lut_adj_427 (.A(\hidden_outputs[1] [10]), .B(n22568), .C(float_alu_c[10]), 
         .D(n70789), .Z(n22569)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_427.init = 16'hc088;
    LUT4 i2_4_lut_adj_428 (.A(n22569), .B(n10_adj_227), .C(\hidden_outputs[1] [10]), 
         .D(n2022[17]), .Z(n62855)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_428.init = 16'hfeee;
    LUT4 i1_4_lut_adj_429 (.A(\hidden_outputs[1] [9]), .B(n22568), .C(float_alu_c[9]), 
         .D(n70789), .Z(n22622)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_429.init = 16'hc088;
    LUT4 i2_4_lut_adj_430 (.A(n10_adj_228), .B(n22622), .C(\hidden_outputs[1] [9]), 
         .D(n2022[17]), .Z(n62907)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_430.init = 16'hfeee;
    LUT4 i1_4_lut_adj_431 (.A(\hidden_outputs[1] [8]), .B(n22568), .C(float_alu_c[8]), 
         .D(n70789), .Z(n22557)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_431.init = 16'hc088;
    LUT4 i1_4_lut_adj_432 (.A(n10_adj_229), .B(\hidden_outputs[1] [8]), 
         .C(n22557), .D(n2022[17]), .Z(n66542)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_432.init = 16'hfefa;
    FD1P3IX n_4659__i21 (.D(n134_adj_403[21]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[21]));
    defparam n_4659__i21.GSR = "DISABLED";
    FD1P3IX n_4659__i20 (.D(n134_adj_403[20]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[20]));
    defparam n_4659__i20.GSR = "DISABLED";
    FD1P3IX n_4659__i19 (.D(n134_adj_403[19]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[19]));
    defparam n_4659__i19.GSR = "DISABLED";
    FD1P3IX n_4659__i18 (.D(n134_adj_403[18]), .SP(n70697), .CD(n24288), 
            .CK(clock), .Q(n[18]));
    defparam n_4659__i18.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_433 (.A(\hidden_outputs[1] [7]), .B(n22568), .C(float_alu_c[7]), 
         .D(n70789), .Z(n23294)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_433.init = 16'hc088;
    PFUMX i54613 (.BLUT(n67522), .ALUT(n67523), .C0(n[1]), .Z(n67524));
    LUT4 i1_4_lut_adj_434 (.A(n10_adj_230), .B(\hidden_outputs[1] [7]), 
         .C(n23294), .D(n2022[17]), .Z(n66540)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_434.init = 16'hfefa;
    LUT4 i1_4_lut_adj_435 (.A(\hidden_outputs[1] [6]), .B(n22568), .C(float_alu_c[6]), 
         .D(n70789), .Z(n22628)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_435.init = 16'hc088;
    PFUMX i54616 (.BLUT(n67525), .ALUT(n67526), .C0(n[1]), .Z(n67527));
    LUT4 i2_4_lut_adj_436 (.A(n10_adj_231), .B(n22628), .C(\hidden_outputs[1] [6]), 
         .D(n2022[17]), .Z(n62909)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_436.init = 16'hfeee;
    LUT4 i1_4_lut_adj_437 (.A(\hidden_outputs[1] [5]), .B(n22568), .C(float_alu_c[5]), 
         .D(n70789), .Z(n23288)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_437.init = 16'hc088;
    LUT4 i2_4_lut_adj_438 (.A(n23288), .B(n10_adj_232), .C(\hidden_outputs[1] [5]), 
         .D(n2022[17]), .Z(n63076)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_438.init = 16'hfeee;
    LUT4 i1_4_lut_adj_439 (.A(\hidden_outputs[1] [4]), .B(n22568), .C(float_alu_c[4]), 
         .D(n70789), .Z(n22631)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_439.init = 16'hc088;
    LUT4 i1_4_lut_adj_440 (.A(n10_adj_233), .B(n22631), .C(\hidden_outputs[1] [4]), 
         .D(n2022[17]), .Z(n66514)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_440.init = 16'hfeee;
    LUT4 i1_4_lut_adj_441 (.A(\hidden_outputs[1] [3]), .B(n22568), .C(float_alu_c[3]), 
         .D(n70789), .Z(n23279)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_441.init = 16'hc088;
    LUT4 i1_4_lut_adj_442 (.A(n10_adj_234), .B(\hidden_outputs[1] [3]), 
         .C(n23279), .D(n2022[17]), .Z(n66278)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_442.init = 16'hfefa;
    LUT4 i1_4_lut_adj_443 (.A(\hidden_outputs[1] [2]), .B(n22568), .C(float_alu_c[2]), 
         .D(n70789), .Z(n22634)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_443.init = 16'hc088;
    LUT4 i2_4_lut_adj_444 (.A(n10_adj_235), .B(n22634), .C(\hidden_outputs[1] [2]), 
         .D(n2022[17]), .Z(n62912)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_444.init = 16'hfeee;
    LUT4 i1_4_lut_adj_445 (.A(\hidden_outputs[1] [1]), .B(n22568), .C(float_alu_c[1]), 
         .D(n70789), .Z(n23276)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_445.init = 16'hc088;
    FD1P3IX counter_4663_4767__i1 (.D(n54[0]), .SP(n4613), .CD(n34857), 
            .CK(clock), .Q(counter[0]));
    defparam counter_4663_4767__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_446 (.A(n10_adj_236), .B(\hidden_outputs[1] [1]), 
         .C(n23276), .D(n2022[17]), .Z(n66284)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_446.init = 16'hfefa;
    LUT4 select_454_Select_31_i10_2_lut (.A(sram_output_B[31]), .B(n2022[9]), 
         .Z(n10_adj_182)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_31_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_447 (.A(\hidden_outputs[0] [31]), .B(n22568), .C(float_alu_c[31]), 
         .D(n70791), .Z(n23249)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_447.init = 16'h88c0;
    LUT4 i2_4_lut_adj_448 (.A(n23249), .B(n10_adj_182), .C(n1586), .D(n2022[17]), 
         .Z(n63060)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_448.init = 16'hfeee;
    LUT4 select_454_Select_30_i10_2_lut (.A(sram_output_B[30]), .B(n2022[9]), 
         .Z(n10_adj_183)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_30_i10_2_lut.init = 16'h8888;
    FD1P3IX i_4655__i0 (.D(n134_adj_409[0]), .SP(n70695), .CD(n23968), 
            .CK(clock), .Q(i[0]));
    defparam i_4655__i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_449 (.A(\hidden_outputs[0] [30]), .B(n22568), .C(float_alu_c[30]), 
         .D(n70791), .Z(n22560)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_449.init = 16'h88c0;
    LUT4 i1_4_lut_adj_450 (.A(n10_adj_183), .B(n22560), .C(\hidden_outputs[0] [30]), 
         .D(n2022[17]), .Z(n66538)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_450.init = 16'hfeee;
    LUT4 select_454_Select_29_i10_2_lut (.A(sram_output_B[29]), .B(n2022[9]), 
         .Z(n10_adj_185)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_29_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_451 (.A(\hidden_outputs[0] [29]), .B(n22568), .C(float_alu_c[29]), 
         .D(n70791), .Z(n23219)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_451.init = 16'h88c0;
    LUT4 i2_4_lut_adj_452 (.A(n23219), .B(n10_adj_185), .C(\hidden_outputs[0] [29]), 
         .D(n2022[17]), .Z(n63052)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_452.init = 16'hfeee;
    LUT4 select_454_Select_28_i10_2_lut (.A(sram_output_B[28]), .B(n2022[9]), 
         .Z(n10_adj_186)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_28_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_453 (.A(\hidden_outputs[0] [28]), .B(n22568), .C(float_alu_c[28]), 
         .D(n70791), .Z(n23213)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_453.init = 16'h88c0;
    LUT4 i2_4_lut_adj_454 (.A(n23213), .B(n10_adj_186), .C(\hidden_outputs[0] [28]), 
         .D(n2022[17]), .Z(n63095)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_454.init = 16'hfeee;
    LUT4 select_454_Select_27_i10_2_lut (.A(sram_output_B[27]), .B(n2022[9]), 
         .Z(n10_adj_187)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_27_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_455 (.A(\hidden_outputs[0] [27]), .B(n22568), .C(float_alu_c[27]), 
         .D(n70791), .Z(n23177)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_455.init = 16'h88c0;
    LUT4 i1_4_lut_adj_456 (.A(n10_adj_187), .B(\hidden_outputs[0] [27]), 
         .C(n23177), .D(n2022[17]), .Z(n66312)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_456.init = 16'hfefa;
    LUT4 select_454_Select_26_i10_2_lut (.A(sram_output_B[26]), .B(n2022[9]), 
         .Z(n10_adj_188)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_26_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_457 (.A(\hidden_outputs[0] [26]), .B(n22568), .C(float_alu_c[26]), 
         .D(n70791), .Z(n23489)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_457.init = 16'h88c0;
    PFUMX i54619 (.BLUT(n67528), .ALUT(n67529), .C0(n[1]), .Z(n67530));
    LUT4 i1_4_lut_adj_458 (.A(n10_adj_188), .B(\hidden_outputs[0] [26]), 
         .C(n23489), .D(n2022[17]), .Z(n66346)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_458.init = 16'hfefa;
    LUT4 select_454_Select_25_i10_2_lut (.A(sram_output_B[25]), .B(n2022[9]), 
         .Z(n10_adj_189)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_25_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_459 (.A(\hidden_outputs[0] [25]), .B(n22568), .C(float_alu_c[25]), 
         .D(n70791), .Z(n22814)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_459.init = 16'h88c0;
    LUT4 i2_4_lut_adj_460 (.A(n10_adj_189), .B(n22814), .C(\hidden_outputs[0] [25]), 
         .D(n2022[17]), .Z(n62971)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_460.init = 16'hfeee;
    LUT4 select_454_Select_24_i10_2_lut (.A(sram_output_B[24]), .B(n2022[9]), 
         .Z(n10_adj_190)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_24_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_461 (.A(\hidden_outputs[0] [24]), .B(n22568), .C(float_alu_c[24]), 
         .D(n70791), .Z(n23171)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_461.init = 16'h88c0;
    LUT4 i2_4_lut_adj_462 (.A(n23171), .B(n10_adj_190), .C(\hidden_outputs[0] [24]), 
         .D(n2022[17]), .Z(n63046)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_462.init = 16'hfeee;
    PFUMX i54622 (.BLUT(n67531), .ALUT(n67532), .C0(n[1]), .Z(n67533));
    LUT4 select_454_Select_23_i10_2_lut (.A(sram_output_B[23]), .B(n2022[9]), 
         .Z(n10_adj_191)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_23_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_463 (.A(\hidden_outputs[0] [23]), .B(n22568), .C(float_alu_c[23]), 
         .D(n70791), .Z(n22820)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_463.init = 16'h88c0;
    LUT4 i1_4_lut_adj_464 (.A(n10_adj_191), .B(n22820), .C(\hidden_outputs[0] [23]), 
         .D(n2022[17]), .Z(n66448)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_464.init = 16'hfeee;
    PFUMX i54625 (.BLUT(n67534), .ALUT(n67535), .C0(n[1]), .Z(n67536));
    PFUMX i54628 (.BLUT(n67537), .ALUT(n67538), .C0(n[1]), .Z(n67539));
    LUT4 select_454_Select_22_i10_2_lut (.A(sram_output_B[22]), .B(n2022[9]), 
         .Z(n10_adj_192)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_22_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_465 (.A(\hidden_outputs[0] [22]), .B(n22568), .C(float_alu_c[22]), 
         .D(n70791), .Z(n23168)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_465.init = 16'h88c0;
    PFUMX i54631 (.BLUT(n67540), .ALUT(n67541), .C0(n[1]), .Z(n67542));
    LUT4 i1_4_lut_adj_466 (.A(n10_adj_192), .B(\hidden_outputs[0] [22]), 
         .C(n23168), .D(n2022[17]), .Z(n66402)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_466.init = 16'hfefa;
    LUT4 select_454_Select_21_i10_2_lut (.A(sram_output_B[21]), .B(n2022[9]), 
         .Z(n10_adj_193)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_21_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_467 (.A(\hidden_outputs[0] [21]), .B(n22568), .C(float_alu_c[21]), 
         .D(n70791), .Z(n22829)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_467.init = 16'h88c0;
    LUT4 i2_4_lut_adj_468 (.A(n10_adj_193), .B(n22829), .C(\hidden_outputs[0] [21]), 
         .D(n2022[17]), .Z(n62975)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_468.init = 16'hfeee;
    LUT4 select_454_Select_20_i10_2_lut (.A(sram_output_B[20]), .B(n2022[9]), 
         .Z(n10_adj_194)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_20_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_469 (.A(\hidden_outputs[0] [20]), .B(n22568), .C(float_alu_c[20]), 
         .D(n70791), .Z(n23462)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_469.init = 16'h88c0;
    LUT4 i1_4_lut_adj_470 (.A(n10_adj_194), .B(\hidden_outputs[0] [20]), 
         .C(n23462), .D(n2022[17]), .Z(n66356)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_470.init = 16'hfefa;
    LUT4 select_454_Select_19_i10_2_lut (.A(sram_output_B[19]), .B(n2022[9]), 
         .Z(n10_adj_195)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_19_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_471 (.A(\hidden_outputs[0] [19]), .B(n22568), .C(float_alu_c[19]), 
         .D(n70791), .Z(n23180)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_471.init = 16'h88c0;
    LUT4 i2_4_lut_adj_472 (.A(n23180), .B(n10_adj_195), .C(\hidden_outputs[0] [19]), 
         .D(n2022[17]), .Z(n63049)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_472.init = 16'hfeee;
    LUT4 select_454_Select_18_i10_2_lut (.A(sram_output_B[18]), .B(n2022[9]), 
         .Z(n10_adj_196)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_18_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_473 (.A(\hidden_outputs[0] [18]), .B(n22568), .C(float_alu_c[18]), 
         .D(n70791), .Z(n23456)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_473.init = 16'h88c0;
    LUT4 i2_4_lut_adj_474 (.A(n23456), .B(n10_adj_196), .C(\hidden_outputs[0] [18]), 
         .D(n2022[17]), .Z(n63224)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_474.init = 16'hfeee;
    LUT4 select_454_Select_17_i10_2_lut (.A(sram_output_B[17]), .B(n2022[9]), 
         .Z(n10_adj_199)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_17_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_475 (.A(\hidden_outputs[0] [17]), .B(n22568), .C(float_alu_c[17]), 
         .D(n70791), .Z(n23453)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_475.init = 16'h88c0;
    LUT4 i2_4_lut_adj_476 (.A(n23453), .B(n10_adj_199), .C(\hidden_outputs[0] [17]), 
         .D(n2022[17]), .Z(n63223)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_476.init = 16'hfeee;
    LUT4 select_454_Select_16_i10_2_lut (.A(sram_output_B[16]), .B(n2022[9]), 
         .Z(n10_adj_205)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_16_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_477 (.A(\hidden_outputs[0] [16]), .B(n22568), .C(float_alu_c[16]), 
         .D(n70791), .Z(n22589)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_477.init = 16'h88c0;
    LUT4 i2_4_lut_adj_478 (.A(n10_adj_205), .B(n22589), .C(\hidden_outputs[0] [16]), 
         .D(n2022[17]), .Z(n62875)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_478.init = 16'hfeee;
    LUT4 select_454_Select_15_i10_2_lut (.A(sram_output_B[15]), .B(n2022[9]), 
         .Z(n10_adj_207)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_15_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_479 (.A(\hidden_outputs[0] [15]), .B(n22568), .C(float_alu_c[15]), 
         .D(n70791), .Z(n23399)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_479.init = 16'h88c0;
    LUT4 i1_4_lut_adj_480 (.A(n10_adj_207), .B(\hidden_outputs[0] [15]), 
         .C(n23399), .D(n2022[17]), .Z(n66374)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_480.init = 16'hfefa;
    LUT4 select_450_Select_14_i10_2_lut (.A(sram_output_B[14]), .B(n2022[9]), 
         .Z(n10_adj_222)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_14_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_481 (.A(\hidden_outputs[0] [14]), .B(n22568), .C(float_alu_c[14]), 
         .D(n70791), .Z(n23135)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_481.init = 16'h88c0;
    LUT4 i2_4_lut_adj_482 (.A(n23135), .B(n10_adj_222), .C(\hidden_outputs[0] [14]), 
         .D(n2022[17]), .Z(n63027)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_482.init = 16'hfeee;
    LUT4 select_450_Select_13_i10_2_lut (.A(sram_output_B[13]), .B(n2022[9]), 
         .Z(n10_adj_224)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_13_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_483 (.A(\hidden_outputs[0] [13]), .B(n22568), .C(float_alu_c[13]), 
         .D(n70791), .Z(n23132)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_483.init = 16'h88c0;
    LUT4 i2_4_lut_adj_484 (.A(n23132), .B(n10_adj_224), .C(\hidden_outputs[0] [13]), 
         .D(n2022[17]), .Z(n63024)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_484.init = 16'hfeee;
    LUT4 select_450_Select_12_i10_2_lut (.A(sram_output_B[12]), .B(n2022[9]), 
         .Z(n10_adj_225)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_12_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_485 (.A(\hidden_outputs[0] [12]), .B(n22568), .C(float_alu_c[12]), 
         .D(n70791), .Z(n22592)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_485.init = 16'h88c0;
    LUT4 i1_4_lut_adj_486 (.A(n10_adj_225), .B(n22592), .C(\hidden_outputs[0] [12]), 
         .D(n2022[17]), .Z(n66444)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_486.init = 16'hfeee;
    CCU2D equal_232_32_49661 (.A0(n[7]), .B0(n[6]), .C0(n[5]), .D0(n[4]), 
          .A1(n[4]), .B1(n[3]), .C1(n[2]), .D1(n[1]), .CIN(n60989), 
          .COUT(n60990));
    defparam equal_232_32_49661.INIT0 = 16'h8001;
    defparam equal_232_32_49661.INIT1 = 16'h8001;
    defparam equal_232_32_49661.INJECT1_0 = "YES";
    defparam equal_232_32_49661.INJECT1_1 = "YES";
    LUT4 select_450_Select_11_i10_2_lut (.A(sram_output_B[11]), .B(n2022[9]), 
         .Z(n10_adj_226)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_11_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_487 (.A(\hidden_outputs[0] [11]), .B(n22568), .C(float_alu_c[11]), 
         .D(n70791), .Z(n23411)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_487.init = 16'h88c0;
    LUT4 i2_4_lut_adj_488 (.A(n23411), .B(n10_adj_226), .C(\hidden_outputs[0] [11]), 
         .D(n2022[17]), .Z(n63207)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_488.init = 16'hfeee;
    LUT4 select_450_Select_10_i10_2_lut (.A(sram_output_B[10]), .B(n2022[9]), 
         .Z(n10_adj_227)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_10_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_489 (.A(\hidden_outputs[0] [10]), .B(n22568), .C(float_alu_c[10]), 
         .D(n70791), .Z(n22871)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_489.init = 16'h88c0;
    LUT4 i2_4_lut_adj_490 (.A(n10_adj_227), .B(n22871), .C(\hidden_outputs[0] [10]), 
         .D(n2022[17]), .Z(n62988)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_490.init = 16'hfeee;
    LUT4 select_450_Select_9_i10_2_lut (.A(sram_output_B[9]), .B(n2022[9]), 
         .Z(n10_adj_228)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_9_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_491 (.A(\hidden_outputs[0] [9]), .B(n22568), .C(float_alu_c[9]), 
         .D(n70791), .Z(n22883)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_491.init = 16'h88c0;
    LUT4 i1_4_lut_adj_492 (.A(n10_adj_228), .B(n22883), .C(\hidden_outputs[0] [9]), 
         .D(n2022[17]), .Z(n66426)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_492.init = 16'hfeee;
    LUT4 select_450_Select_8_i10_2_lut (.A(sram_output_B[8]), .B(n2022[9]), 
         .Z(n10_adj_229)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_8_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_493 (.A(\hidden_outputs[0] [8]), .B(n22568), .C(float_alu_c[8]), 
         .D(n70791), .Z(n22880)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_493.init = 16'h88c0;
    LUT4 i1_4_lut_adj_494 (.A(n10_adj_229), .B(n22880), .C(\hidden_outputs[0] [8]), 
         .D(n2022[17]), .Z(n66428)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_494.init = 16'hfeee;
    LUT4 select_450_Select_7_i10_2_lut (.A(sram_output_B[7]), .B(n2022[9]), 
         .Z(n10_adj_230)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_7_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_495 (.A(\hidden_outputs[0] [7]), .B(n22568), .C(float_alu_c[7]), 
         .D(n70791), .Z(n22889)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_495.init = 16'h88c0;
    LUT4 i2_4_lut_adj_496 (.A(n10_adj_230), .B(n22889), .C(\hidden_outputs[0] [7]), 
         .D(n2022[17]), .Z(n63000)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_496.init = 16'hfeee;
    LUT4 select_450_Select_6_i10_2_lut (.A(sram_output_B[6]), .B(n2022[9]), 
         .Z(n10_adj_231)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_6_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_497 (.A(\hidden_outputs[0] [6]), .B(n22568), .C(float_alu_c[6]), 
         .D(n70791), .Z(n22886)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_497.init = 16'h88c0;
    LUT4 i1_4_lut_adj_498 (.A(n10_adj_231), .B(n22886), .C(\hidden_outputs[0] [6]), 
         .D(n2022[17]), .Z(n66422)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_498.init = 16'hfeee;
    LUT4 select_450_Select_5_i10_2_lut (.A(sram_output_B[5]), .B(n2022[9]), 
         .Z(n10_adj_232)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_5_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_499 (.A(\hidden_outputs[0] [5]), .B(n22568), .C(float_alu_c[5]), 
         .D(n70791), .Z(n22892)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_499.init = 16'h88c0;
    LUT4 i1_4_lut_adj_500 (.A(n10_adj_232), .B(n22892), .C(\hidden_outputs[0] [5]), 
         .D(n2022[17]), .Z(n66420)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_500.init = 16'hfeee;
    LUT4 select_450_Select_4_i10_2_lut (.A(sram_output_B[4]), .B(n2022[9]), 
         .Z(n10_adj_233)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_4_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_501 (.A(\hidden_outputs[0] [4]), .B(n22568), .C(float_alu_c[4]), 
         .D(n70791), .Z(n22895)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_501.init = 16'h88c0;
    LUT4 i2_4_lut_adj_502 (.A(n10_adj_233), .B(n22895), .C(\hidden_outputs[0] [4]), 
         .D(n2022[17]), .Z(n63002)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_502.init = 16'hfeee;
    LUT4 select_450_Select_3_i10_2_lut (.A(sram_output_B[3]), .B(n2022[9]), 
         .Z(n10_adj_234)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_450_Select_3_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_503 (.A(\hidden_outputs[0] [3]), .B(n22568), .C(float_alu_c[3]), 
         .D(n70791), .Z(n23129)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_503.init = 16'h88c0;
    LUT4 i1_4_lut_adj_504 (.A(n10_adj_234), .B(\hidden_outputs[0] [3]), 
         .C(n23129), .D(n2022[17]), .Z(n66548)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_504.init = 16'hfefa;
    LUT4 select_454_Select_2_i10_2_lut (.A(sram_output_B[2]), .B(n2022[9]), 
         .Z(n10_adj_235)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_2_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_505 (.A(\hidden_outputs[0] [2]), .B(n22568), .C(float_alu_c[2]), 
         .D(n70791), .Z(n22595)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_505.init = 16'h88c0;
    LUT4 i1_4_lut_adj_506 (.A(n10_adj_235), .B(n22595), .C(\hidden_outputs[0] [2]), 
         .D(n2022[17]), .Z(n66528)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_506.init = 16'hfeee;
    LUT4 i54486_3_lut (.A(\hidden_outputs[2] [14]), .B(\hidden_outputs[3] [14]), 
         .C(h[0]), .Z(n67397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54486_3_lut.init = 16'hcaca;
    LUT4 i54485_3_lut (.A(\hidden_outputs[0] [14]), .B(\hidden_outputs[1] [14]), 
         .C(h[0]), .Z(n67396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54485_3_lut.init = 16'hcaca;
    LUT4 i54483_3_lut (.A(\hidden_outputs[2] [13]), .B(\hidden_outputs[3] [13]), 
         .C(h[0]), .Z(n67394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54483_3_lut.init = 16'hcaca;
    LUT4 i54482_3_lut (.A(\hidden_outputs[0] [13]), .B(\hidden_outputs[1] [13]), 
         .C(h[0]), .Z(n67393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54482_3_lut.init = 16'hcaca;
    LUT4 i54480_3_lut (.A(\hidden_outputs[2] [12]), .B(\hidden_outputs[3] [12]), 
         .C(h[0]), .Z(n67391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54480_3_lut.init = 16'hcaca;
    LUT4 i54479_3_lut (.A(\hidden_outputs[0] [12]), .B(\hidden_outputs[1] [12]), 
         .C(h[0]), .Z(n67390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54479_3_lut.init = 16'hcaca;
    LUT4 i54477_3_lut (.A(\hidden_outputs[2] [11]), .B(\hidden_outputs[3] [11]), 
         .C(h[0]), .Z(n67388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54477_3_lut.init = 16'hcaca;
    LUT4 i54476_3_lut (.A(\hidden_outputs[0] [11]), .B(\hidden_outputs[1] [11]), 
         .C(h[0]), .Z(n67387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54476_3_lut.init = 16'hcaca;
    LUT4 i54474_3_lut (.A(\hidden_outputs[2] [10]), .B(\hidden_outputs[3] [10]), 
         .C(h[0]), .Z(n67385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54474_3_lut.init = 16'hcaca;
    LUT4 i54473_3_lut (.A(\hidden_outputs[0] [10]), .B(\hidden_outputs[1] [10]), 
         .C(h[0]), .Z(n67384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54473_3_lut.init = 16'hcaca;
    LUT4 i54471_3_lut (.A(\hidden_outputs[2] [9]), .B(\hidden_outputs[3] [9]), 
         .C(h[0]), .Z(n67382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54471_3_lut.init = 16'hcaca;
    LUT4 i54470_3_lut (.A(\hidden_outputs[0] [9]), .B(\hidden_outputs[1] [9]), 
         .C(h[0]), .Z(n67381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54470_3_lut.init = 16'hcaca;
    LUT4 i54468_3_lut (.A(\hidden_outputs[2] [8]), .B(\hidden_outputs[3] [8]), 
         .C(h[0]), .Z(n67379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54468_3_lut.init = 16'hcaca;
    LUT4 i54467_3_lut (.A(\hidden_outputs[0] [8]), .B(\hidden_outputs[1] [8]), 
         .C(h[0]), .Z(n67378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54467_3_lut.init = 16'hcaca;
    LUT4 i54465_3_lut (.A(\hidden_outputs[2] [7]), .B(\hidden_outputs[3] [7]), 
         .C(h[0]), .Z(n67376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54465_3_lut.init = 16'hcaca;
    LUT4 i54464_3_lut (.A(\hidden_outputs[0] [7]), .B(\hidden_outputs[1] [7]), 
         .C(h[0]), .Z(n67375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54464_3_lut.init = 16'hcaca;
    LUT4 i54462_3_lut (.A(\hidden_outputs[2] [6]), .B(\hidden_outputs[3] [6]), 
         .C(h[0]), .Z(n67373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54462_3_lut.init = 16'hcaca;
    LUT4 i54461_3_lut (.A(\hidden_outputs[0] [6]), .B(\hidden_outputs[1] [6]), 
         .C(h[0]), .Z(n67372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54461_3_lut.init = 16'hcaca;
    LUT4 i54459_3_lut (.A(\hidden_outputs[2] [5]), .B(\hidden_outputs[3] [5]), 
         .C(h[0]), .Z(n67370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54459_3_lut.init = 16'hcaca;
    LUT4 i54458_3_lut (.A(\hidden_outputs[0] [5]), .B(\hidden_outputs[1] [5]), 
         .C(h[0]), .Z(n67369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54458_3_lut.init = 16'hcaca;
    LUT4 i54456_3_lut (.A(\hidden_outputs[2] [4]), .B(\hidden_outputs[3] [4]), 
         .C(h[0]), .Z(n67367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54456_3_lut.init = 16'hcaca;
    LUT4 i54455_3_lut (.A(\hidden_outputs[0] [4]), .B(\hidden_outputs[1] [4]), 
         .C(h[0]), .Z(n67366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54455_3_lut.init = 16'hcaca;
    LUT4 i54453_3_lut (.A(\hidden_outputs[2] [3]), .B(\hidden_outputs[3] [3]), 
         .C(h[0]), .Z(n67364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54453_3_lut.init = 16'hcaca;
    LUT4 i54452_3_lut (.A(\hidden_outputs[0] [3]), .B(\hidden_outputs[1] [3]), 
         .C(h[0]), .Z(n67363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54452_3_lut.init = 16'hcaca;
    LUT4 i54450_3_lut (.A(\hidden_outputs[2] [2]), .B(\hidden_outputs[3] [2]), 
         .C(h[0]), .Z(n67361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54450_3_lut.init = 16'hcaca;
    LUT4 i54449_3_lut (.A(\hidden_outputs[0] [2]), .B(\hidden_outputs[1] [2]), 
         .C(h[0]), .Z(n67360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54449_3_lut.init = 16'hcaca;
    LUT4 i54447_3_lut (.A(\hidden_outputs[2] [1]), .B(\hidden_outputs[3] [1]), 
         .C(h[0]), .Z(n67358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54447_3_lut.init = 16'hcaca;
    LUT4 i54446_3_lut (.A(\hidden_outputs[0] [1]), .B(\hidden_outputs[1] [1]), 
         .C(h[0]), .Z(n67357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54446_3_lut.init = 16'hcaca;
    LUT4 i54444_3_lut (.A(\temp_outputs[2] [1]), .B(\temp_outputs[3] [1]), 
         .C(i[0]), .Z(n67355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54444_3_lut.init = 16'hcaca;
    LUT4 i54443_3_lut (.A(\temp_outputs[0] [1]), .B(\temp_outputs[1] [1]), 
         .C(i[0]), .Z(n67354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54443_3_lut.init = 16'hcaca;
    LUT4 i54441_3_lut (.A(\temp_outputs[2] [2]), .B(\temp_outputs[3] [2]), 
         .C(i[0]), .Z(n67352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54441_3_lut.init = 16'hcaca;
    LUT4 i54440_3_lut (.A(\temp_outputs[0] [2]), .B(\temp_outputs[1] [2]), 
         .C(i[0]), .Z(n67351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54440_3_lut.init = 16'hcaca;
    LUT4 mux_141_Mux_24_i7_4_lut (.A(n67428), .B(\hidden_outputs[4] [24]), 
         .C(h[2]), .D(n70861), .Z(n2448[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_24_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_24_i1_3_lut (.A(\mlp_outputs[0] [24]), .B(\mlp_outputs[1] [24]), 
         .C(o[0]), .Z(n4478[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_24_i1_3_lut.init = 16'hcaca;
    LUT4 mux_75_Mux_24_i7_4_lut (.A(n67290), .B(\temp_outputs[4] [24]), 
         .C(i[2]), .D(n17802), .Z(n1028[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_24_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i25_3_lut (.A(n1028[24]), .B(n1027[24]), .C(n70712), .Z(n1061[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i25_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_507 (.A(n2448[24]), .B(e[24]), .C(n70864), .D(n2022[15]), 
         .Z(n8_adj_349)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_507.init = 16'heca0;
    LUT4 select_460_Select_24_i38_2_lut (.A(f[24]), .B(n2022[37]), .Z(n38_adj_350)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_24_i38_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_508 (.A(n17650), .B(n8_adj_349), .C(n1061[24]), 
         .D(n2022[13]), .Z(n10_adj_351)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_508.init = 16'hfeee;
    LUT4 mux_220_Mux_24_i7_4_lut (.A(n67521), .B(\hidden_outputs[4] [24]), 
         .C(n[2]), .D(n70842), .Z(n3742[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_24_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_509 (.A(n3742[24]), .B(n10_adj_351), .C(n38_adj_350), 
         .D(n2022[35]), .Z(n63254)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_509.init = 16'hfefc;
    LUT4 mux_75_Mux_28_i7_4_lut (.A(n67278), .B(\temp_outputs[4] [28]), 
         .C(i[2]), .D(n17802), .Z(n1028[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_75_Mux_28_i7_4_lut.init = 16'h0aca;
    LUT4 mux_76_i29_3_lut (.A(n1028[28]), .B(n1027[28]), .C(n70712), .Z(n1061[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mux_76_i29_3_lut.init = 16'hacac;
    LUT4 i2_4_lut_adj_510 (.A(n2448[28]), .B(e[28]), .C(n70864), .D(n2022[15]), 
         .Z(n8_adj_352)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_510.init = 16'heca0;
    LUT4 select_460_Select_28_i38_2_lut (.A(f[28]), .B(n2022[37]), .Z(n38_adj_353)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_460_Select_28_i38_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_511 (.A(n17704), .B(n8_adj_352), .C(n1061[28]), 
         .D(n2022[13]), .Z(n10_adj_354)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i4_4_lut_adj_511.init = 16'hfeee;
    LUT4 mux_220_Mux_28_i7_4_lut (.A(n67533), .B(\hidden_outputs[4] [28]), 
         .C(n[2]), .D(n70842), .Z(n3742[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_220_Mux_28_i7_4_lut.init = 16'h0aca;
    LUT4 i5_4_lut_adj_512 (.A(n3742[28]), .B(n10_adj_354), .C(n38_adj_353), 
         .D(n2022[35]), .Z(n63159)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_512.init = 16'hfefc;
    LUT4 i2_4_lut_adj_513 (.A(n70822), .B(n70858), .C(n70736), .D(n70857), 
         .Z(n63295)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i2_4_lut_adj_513.init = 16'ha888;
    LUT4 i54438_3_lut (.A(\temp_outputs[2] [3]), .B(\temp_outputs[3] [3]), 
         .C(i[0]), .Z(n67349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54438_3_lut.init = 16'hcaca;
    LUT4 i54437_3_lut (.A(\temp_outputs[0] [3]), .B(\temp_outputs[1] [3]), 
         .C(i[0]), .Z(n67348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54437_3_lut.init = 16'hcaca;
    LUT4 i54435_3_lut (.A(\temp_outputs[2] [4]), .B(\temp_outputs[3] [4]), 
         .C(i[0]), .Z(n67346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54435_3_lut.init = 16'hcaca;
    LUT4 i54434_3_lut (.A(\temp_outputs[0] [4]), .B(\temp_outputs[1] [4]), 
         .C(i[0]), .Z(n67345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54434_3_lut.init = 16'hcaca;
    LUT4 i54432_3_lut (.A(\temp_outputs[2] [5]), .B(\temp_outputs[3] [5]), 
         .C(i[0]), .Z(n67343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54432_3_lut.init = 16'hcaca;
    LUT4 i54431_3_lut (.A(\temp_outputs[0] [5]), .B(\temp_outputs[1] [5]), 
         .C(i[0]), .Z(n67342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54431_3_lut.init = 16'hcaca;
    LUT4 i54429_3_lut (.A(\temp_outputs[2] [6]), .B(\temp_outputs[3] [6]), 
         .C(i[0]), .Z(n67340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54429_3_lut.init = 16'hcaca;
    LUT4 i54428_3_lut (.A(\temp_outputs[0] [6]), .B(\temp_outputs[1] [6]), 
         .C(i[0]), .Z(n67339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54428_3_lut.init = 16'hcaca;
    LUT4 i54426_3_lut (.A(\temp_outputs[2] [7]), .B(\temp_outputs[3] [7]), 
         .C(i[0]), .Z(n67337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54426_3_lut.init = 16'hcaca;
    LUT4 i54425_3_lut (.A(\temp_outputs[0] [7]), .B(\temp_outputs[1] [7]), 
         .C(i[0]), .Z(n67336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54425_3_lut.init = 16'hcaca;
    LUT4 i54423_3_lut (.A(\temp_outputs[2] [8]), .B(\temp_outputs[3] [8]), 
         .C(i[0]), .Z(n67334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54423_3_lut.init = 16'hcaca;
    LUT4 i54422_3_lut (.A(\temp_outputs[0] [8]), .B(\temp_outputs[1] [8]), 
         .C(i[0]), .Z(n67333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54422_3_lut.init = 16'hcaca;
    LUT4 i54420_3_lut (.A(\temp_outputs[2] [9]), .B(\temp_outputs[3] [9]), 
         .C(i[0]), .Z(n67331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54420_3_lut.init = 16'hcaca;
    LUT4 i54419_3_lut (.A(\temp_outputs[0] [9]), .B(\temp_outputs[1] [9]), 
         .C(i[0]), .Z(n67330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54419_3_lut.init = 16'hcaca;
    LUT4 i54417_3_lut (.A(\temp_outputs[2] [10]), .B(\temp_outputs[3] [10]), 
         .C(i[0]), .Z(n67328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54417_3_lut.init = 16'hcaca;
    LUT4 i54416_3_lut (.A(\temp_outputs[0] [10]), .B(\temp_outputs[1] [10]), 
         .C(i[0]), .Z(n67327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54416_3_lut.init = 16'hcaca;
    LUT4 i54414_3_lut (.A(\temp_outputs[2] [11]), .B(\temp_outputs[3] [11]), 
         .C(i[0]), .Z(n67325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54414_3_lut.init = 16'hcaca;
    LUT4 i54413_3_lut (.A(\temp_outputs[0] [11]), .B(\temp_outputs[1] [11]), 
         .C(i[0]), .Z(n67324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54413_3_lut.init = 16'hcaca;
    LUT4 i54411_3_lut (.A(\temp_outputs[2] [12]), .B(\temp_outputs[3] [12]), 
         .C(i[0]), .Z(n67322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54411_3_lut.init = 16'hcaca;
    LUT4 i54410_3_lut (.A(\temp_outputs[0] [12]), .B(\temp_outputs[1] [12]), 
         .C(i[0]), .Z(n67321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54410_3_lut.init = 16'hcaca;
    LUT4 i54408_3_lut (.A(\temp_outputs[2] [13]), .B(\temp_outputs[3] [13]), 
         .C(i[0]), .Z(n67319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54408_3_lut.init = 16'hcaca;
    LUT4 i54407_3_lut (.A(\temp_outputs[0] [13]), .B(\temp_outputs[1] [13]), 
         .C(i[0]), .Z(n67318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54407_3_lut.init = 16'hcaca;
    LUT4 i54405_3_lut (.A(\temp_outputs[2] [14]), .B(\temp_outputs[3] [14]), 
         .C(i[0]), .Z(n67316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54405_3_lut.init = 16'hcaca;
    LUT4 i54404_3_lut (.A(\temp_outputs[0] [14]), .B(\temp_outputs[1] [14]), 
         .C(i[0]), .Z(n67315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54404_3_lut.init = 16'hcaca;
    LUT4 i54402_3_lut (.A(\temp_outputs[2] [15]), .B(\temp_outputs[3] [15]), 
         .C(i[0]), .Z(n67313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54402_3_lut.init = 16'hcaca;
    LUT4 i54401_3_lut (.A(\temp_outputs[0] [15]), .B(\temp_outputs[1] [15]), 
         .C(i[0]), .Z(n67312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54401_3_lut.init = 16'hcaca;
    CCU2D equal_232_30 (.A0(n[13]), .B0(n[12]), .C0(n[11]), .D0(n[10]), 
          .A1(n[10]), .B1(n[9]), .C1(n[8]), .D1(n[7]), .CIN(n60988), 
          .COUT(n60989));
    defparam equal_232_30.INIT0 = 16'h8001;
    defparam equal_232_30.INIT1 = 16'h8001;
    defparam equal_232_30.INJECT1_0 = "YES";
    defparam equal_232_30.INJECT1_1 = "YES";
    LUT4 i54399_3_lut (.A(\temp_outputs[2] [16]), .B(\temp_outputs[3] [16]), 
         .C(i[0]), .Z(n67310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54399_3_lut.init = 16'hcaca;
    LUT4 i54398_3_lut (.A(\temp_outputs[0] [16]), .B(\temp_outputs[1] [16]), 
         .C(i[0]), .Z(n67309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54398_3_lut.init = 16'hcaca;
    LUT4 i54396_3_lut (.A(\temp_outputs[2] [17]), .B(\temp_outputs[3] [17]), 
         .C(i[0]), .Z(n67307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54396_3_lut.init = 16'hcaca;
    CCU2D equal_232_28 (.A0(n[19]), .B0(n[18]), .C0(n[17]), .D0(n[16]), 
          .A1(n[16]), .B1(n[15]), .C1(n[14]), .D1(n[13]), .CIN(n60987), 
          .COUT(n60988));
    defparam equal_232_28.INIT0 = 16'h8001;
    defparam equal_232_28.INIT1 = 16'h8001;
    defparam equal_232_28.INJECT1_0 = "YES";
    defparam equal_232_28.INJECT1_1 = "YES";
    LUT4 i54395_3_lut (.A(\temp_outputs[0] [17]), .B(\temp_outputs[1] [17]), 
         .C(i[0]), .Z(n67306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54395_3_lut.init = 16'hcaca;
    LUT4 i54393_3_lut (.A(\temp_outputs[2] [18]), .B(\temp_outputs[3] [18]), 
         .C(i[0]), .Z(n67304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54393_3_lut.init = 16'hcaca;
    LUT4 i54392_3_lut (.A(\temp_outputs[0] [18]), .B(\temp_outputs[1] [18]), 
         .C(i[0]), .Z(n67303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54392_3_lut.init = 16'hcaca;
    LUT4 i54390_3_lut (.A(\temp_outputs[2] [19]), .B(\temp_outputs[3] [19]), 
         .C(i[0]), .Z(n67301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54390_3_lut.init = 16'hcaca;
    LUT4 i54389_3_lut (.A(\temp_outputs[0] [19]), .B(\temp_outputs[1] [19]), 
         .C(i[0]), .Z(n67300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54389_3_lut.init = 16'hcaca;
    LUT4 i54387_3_lut (.A(\temp_outputs[2] [21]), .B(\temp_outputs[3] [21]), 
         .C(i[0]), .Z(n67298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54387_3_lut.init = 16'hcaca;
    LUT4 i54386_3_lut (.A(\temp_outputs[0] [21]), .B(\temp_outputs[1] [21]), 
         .C(i[0]), .Z(n67297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54386_3_lut.init = 16'hcaca;
    LUT4 select_454_Select_1_i10_2_lut (.A(sram_output_B[1]), .B(n2022[9]), 
         .Z(n10_adj_236)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_454_Select_1_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_514 (.A(\hidden_outputs[0] [1]), .B(n22568), .C(float_alu_c[1]), 
         .D(n70791), .Z(n22865)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_514.init = 16'h88c0;
    LUT4 i2_4_lut_adj_515 (.A(n22865), .B(n10_adj_236), .C(\hidden_outputs[0] [1]), 
         .D(n2022[17]), .Z(n62897)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_515.init = 16'hfeee;
    LUT4 i54384_3_lut (.A(\temp_outputs[2] [22]), .B(\temp_outputs[3] [22]), 
         .C(i[0]), .Z(n67295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54384_3_lut.init = 16'hcaca;
    LUT4 i54383_3_lut (.A(\temp_outputs[0] [22]), .B(\temp_outputs[1] [22]), 
         .C(i[0]), .Z(n67294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54383_3_lut.init = 16'hcaca;
    CCU2D equal_232_26 (.A0(n[25]), .B0(n[24]), .C0(n[23]), .D0(n[22]), 
          .A1(n[22]), .B1(n[21]), .C1(n[20]), .D1(n[19]), .CIN(n60986), 
          .COUT(n60987));
    defparam equal_232_26.INIT0 = 16'h8001;
    defparam equal_232_26.INIT1 = 16'h8001;
    defparam equal_232_26.INJECT1_0 = "YES";
    defparam equal_232_26.INJECT1_1 = "YES";
    LUT4 i54381_3_lut (.A(\temp_outputs[2] [23]), .B(\temp_outputs[3] [23]), 
         .C(i[0]), .Z(n67292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54381_3_lut.init = 16'hcaca;
    LUT4 i54380_3_lut (.A(\temp_outputs[0] [23]), .B(\temp_outputs[1] [23]), 
         .C(i[0]), .Z(n67291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54380_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_516 (.A(n11102[1]), .B(n61278[1]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_355)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_516.init = 16'heca0;
    LUT4 i2_4_lut_adj_517 (.A(n61250[1]), .B(addr[1]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_356)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_517.init = 16'heca0;
    LUT4 i4_4_lut_adj_518 (.A(n7_adj_356), .B(n61312[1]), .C(n6_adj_355), 
         .D(n2022[32]), .Z(n63018)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_518.init = 16'hfefa;
    LUT4 i1_4_lut_adj_519 (.A(n11102[2]), .B(n61278[2]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_357)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_519.init = 16'heca0;
    LUT4 i2_4_lut_adj_520 (.A(n61250[2]), .B(addr[2]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_358)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_520.init = 16'heca0;
    LUT4 i4_4_lut_adj_521 (.A(n7_adj_358), .B(n61312[2]), .C(n6_adj_357), 
         .D(n2022[32]), .Z(n63135)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_521.init = 16'hfefa;
    LUT4 i1_4_lut_adj_522 (.A(n11102[3]), .B(n61278[3]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_359)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_522.init = 16'heca0;
    LUT4 i2_4_lut_adj_523 (.A(n61250[3]), .B(addr[3]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_360)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_523.init = 16'heca0;
    LUT4 i4_4_lut_adj_524 (.A(n7_adj_360), .B(n61312[3]), .C(n6_adj_359), 
         .D(n2022[32]), .Z(n63138)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_524.init = 16'hfefa;
    LUT4 i1_4_lut_adj_525 (.A(n11102[4]), .B(n61278[4]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_361)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_525.init = 16'heca0;
    LUT4 i2_4_lut_adj_526 (.A(n61250[4]), .B(addr[4]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_362)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_526.init = 16'heca0;
    LUT4 i4_4_lut_adj_527 (.A(n7_adj_362), .B(n61312[4]), .C(n6_adj_361), 
         .D(n2022[32]), .Z(n63238)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_527.init = 16'hfefa;
    LUT4 i1_2_lut_adj_528 (.A(n2036), .B(mlp_mode), .Z(n2242)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_528.init = 16'h8888;
    LUT4 i2_4_lut_adj_529 (.A(n2022[27]), .B(n2082), .C(n2664), .D(n35), 
         .Z(n63041)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(D))) */ ;
    defparam i2_4_lut_adj_529.init = 16'hffce;
    LUT4 i1_2_lut_adj_530 (.A(n2022[9]), .B(n70700), .Z(n2251)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_530.init = 16'heeee;
    LUT4 i6_2_lut (.A(i_c[21]), .B(i_c[25]), .Z(n38_adj_363)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(i_c[26]), .B(i_c[31]), .C(i_c[18]), .D(\i[5] ), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i14_2_lut_adj_531 (.A(i[1]), .B(\i[4] ), .Z(n46_adj_364)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14_2_lut_adj_531.init = 16'heeee;
    LUT4 i24_4_lut_adj_532 (.A(i_c[13]), .B(i[10]), .C(i_c[23]), .D(i_c[20]), 
         .Z(n56_adj_365)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut_adj_532.init = 16'hfffe;
    LUT4 i10_2_lut_adj_533 (.A(i_c[16]), .B(i_c[14]), .Z(n42_adj_366)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i10_2_lut_adj_533.init = 16'heeee;
    LUT4 i22_4_lut_adj_534 (.A(i_c[19]), .B(i_c[27]), .C(i_c[22]), .D(\i[12] ), 
         .Z(n54_adj_367)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut_adj_534.init = 16'hfffe;
    LUT4 i28_4_lut_adj_535 (.A(i_c[17]), .B(n56_adj_365), .C(n46_adj_364), 
         .D(i_c[24]), .Z(n60_adj_368)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i28_4_lut_adj_535.init = 16'hfffe;
    LUT4 i9_2_lut_adj_536 (.A(i[2]), .B(\i[8] ), .Z(n41_adj_369)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i9_2_lut_adj_536.init = 16'hdddd;
    LUT4 i18_4_lut_adj_537 (.A(\i[7] ), .B(\i[3] ), .C(i_c[15]), .D(i_c[29]), 
         .Z(n50_adj_370)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut_adj_537.init = 16'hfffe;
    LUT4 i26_4_lut_adj_538 (.A(i[0]), .B(n52), .C(n38_adj_363), .D(\i[6] ), 
         .Z(n58_adj_371)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut_adj_538.init = 16'hfffe;
    LUT4 i30_4_lut_adj_539 (.A(n41_adj_369), .B(n60_adj_368), .C(n54_adj_367), 
         .D(n42_adj_366), .Z(n62_adj_372)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut_adj_539.init = 16'hfffe;
    LUT4 i17_4_lut_adj_540 (.A(\i[11] ), .B(\i[9] ), .C(i_c[30]), .D(i_c[28]), 
         .Z(n49_adj_373)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_540.init = 16'hfffe;
    LUT4 i31_4_lut_adj_541 (.A(n49_adj_373), .B(n62_adj_372), .C(n58_adj_371), 
         .D(n50_adj_370), .Z(n23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31_4_lut_adj_541.init = 16'hfffe;
    CCU2D equal_232_24 (.A0(n[31]), .B0(n[30]), .C0(n[29]), .D0(n[28]), 
          .A1(n[28]), .B1(n[27]), .C1(n[26]), .D1(n[25]), .CIN(n60985), 
          .COUT(n60986));
    defparam equal_232_24.INIT0 = 16'h8001;
    defparam equal_232_24.INIT1 = 16'h8001;
    defparam equal_232_24.INJECT1_0 = "YES";
    defparam equal_232_24.INJECT1_1 = "YES";
    LUT4 i1_4_lut_adj_542 (.A(n11102[5]), .B(n61278[5]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_374)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_542.init = 16'heca0;
    LUT4 i2_4_lut_adj_543 (.A(n61250[5]), .B(addr[5]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_375)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_543.init = 16'heca0;
    LUT4 i4_4_lut_adj_544 (.A(n7_adj_375), .B(n61312[5]), .C(n6_adj_374), 
         .D(n2022[32]), .Z(n63255)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_544.init = 16'hfefa;
    LUT4 i1_2_lut_adj_545 (.A(n2022[38]), .B(n3922), .Z(n2284)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_545.init = 16'h8888;
    LUT4 i53932_2_lut (.A(o[15]), .B(o[26]), .Z(n66837)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53932_2_lut.init = 16'heeee;
    LUT4 i54066_4_lut (.A(o[14]), .B(o[16]), .C(o[18]), .D(o[6]), .Z(n66975)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54066_4_lut.init = 16'hfffe;
    LUT4 i53940_2_lut (.A(o[30]), .B(o[27]), .Z(n66845)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53940_2_lut.init = 16'heeee;
    LUT4 i54070_4_lut (.A(o[21]), .B(o[31]), .C(o[12]), .D(o[24]), .Z(n66979)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54070_4_lut.init = 16'hfffe;
    LUT4 i54102_4_lut (.A(o[23]), .B(n66975), .C(n66837), .D(o[7]), 
         .Z(n67013)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54102_4_lut.init = 16'hfffe;
    LUT4 i53942_2_lut (.A(o[20]), .B(o[13]), .Z(n66847)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53942_2_lut.init = 16'heeee;
    LUT4 i54078_4_lut (.A(o[1]), .B(o[29]), .C(o[2]), .D(o[8]), .Z(n66987)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54078_4_lut.init = 16'hfffe;
    LUT4 i54074_4_lut (.A(o[22]), .B(o[11]), .C(o[28]), .D(o[25]), .Z(n66983)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54074_4_lut.init = 16'hfffe;
    LUT4 i54076_4_lut (.A(o[19]), .B(o[4]), .C(o[3]), .D(o[10]), .Z(n66985)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54076_4_lut.init = 16'hfffe;
    LUT4 i54118_4_lut (.A(n66847), .B(n67013), .C(n66979), .D(n66845), 
         .Z(n67029)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54118_4_lut.init = 16'hfffe;
    LUT4 i54108_4_lut (.A(o[9]), .B(n66987), .C(o[5]), .D(o[17]), .Z(n67019)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54108_4_lut.init = 16'hfffe;
    LUT4 i54126_4_lut (.A(n67019), .B(n67029), .C(n66985), .D(n66983), 
         .Z(n67037)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i54126_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_adj_546 (.A(n67037), .B(o[0]), .C(n2022[49]), .Z(n63590)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_3_lut_adj_546.init = 16'h4040;
    LUT4 i1_4_lut_adj_547 (.A(n70848), .B(n63590), .C(n2022[3]), .D(n65), 
         .Z(n66556)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i1_4_lut_adj_547.init = 16'heefe;
    LUT4 i1_4_lut_adj_548 (.A(n11102[6]), .B(n61278[6]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_376)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_548.init = 16'heca0;
    LUT4 i2_4_lut_adj_549 (.A(n61250[6]), .B(addr[6]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_377)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_549.init = 16'heca0;
    LUT4 i4_4_lut_adj_550 (.A(n7_adj_377), .B(n61312[6]), .C(n6_adj_376), 
         .D(n2022[32]), .Z(n63167)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_550.init = 16'hfefa;
    LUT4 i1_4_lut_adj_551 (.A(n11102[7]), .B(n61278[7]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_378)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_551.init = 16'heca0;
    LUT4 i2_4_lut_adj_552 (.A(n61250[7]), .B(addr[7]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_379)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_552.init = 16'heca0;
    LUT4 i4_4_lut_adj_553 (.A(n7_adj_379), .B(n61312[7]), .C(n6_adj_378), 
         .D(n2022[32]), .Z(n63164)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_553.init = 16'hfefa;
    LUT4 i12330_4_lut (.A(n23680), .B(n2022[27]), .C(n2664), .D(n2022[28]), 
         .Z(n24020)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i12330_4_lut.init = 16'haaa2;
    LUT4 i22_3_lut (.A(n2082), .B(n2664), .C(n2022[27]), .Z(n12_adj_380)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i22_3_lut.init = 16'h3a3a;
    LUT4 i1_4_lut_adj_554 (.A(n12_adj_380), .B(n70822), .C(n70713), .D(n2022[28]), 
         .Z(n23680)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_554.init = 16'hc088;
    LUT4 i1_4_lut_adj_555 (.A(n11102[8]), .B(n61278[8]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_381)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_555.init = 16'heca0;
    LUT4 i2_4_lut_adj_556 (.A(n61250[8]), .B(addr[8]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_382)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_556.init = 16'heca0;
    LUT4 i4_4_lut_adj_557 (.A(n7_adj_382), .B(n61312[8]), .C(n6_adj_381), 
         .D(n2022[32]), .Z(n63163)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_557.init = 16'hfefa;
    LUT4 i1_4_lut_adj_558 (.A(n11102[9]), .B(n61278[9]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_383)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_558.init = 16'heca0;
    LUT4 i2_4_lut_adj_559 (.A(n61250[9]), .B(addr[9]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_384)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_559.init = 16'heca0;
    LUT4 i4_4_lut_adj_560 (.A(n7_adj_384), .B(n61312[9]), .C(n6_adj_383), 
         .D(n2022[32]), .Z(n63158)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_560.init = 16'hfefa;
    LUT4 i11_2_lut (.A(addr[25]), .B(addr[27]), .Z(n40_adj_385)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11_2_lut.init = 16'heeee;
    LUT4 i21_4_lut_adj_561 (.A(addr[28]), .B(addr[23]), .C(addr[2]), .D(addr[24]), 
         .Z(n50_adj_386)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut_adj_561.init = 16'hfffe;
    LUT4 i7_2_lut_adj_562 (.A(addr[9]), .B(addr[12]), .Z(n36_adj_387)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_adj_562.init = 16'heeee;
    LUT4 i19_4_lut_adj_563 (.A(addr[14]), .B(addr[8]), .C(addr[5]), .D(addr[29]), 
         .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut_adj_563.init = 16'hfffe;
    LUT4 i3_2_lut (.A(addr[19]), .B(addr[20]), .Z(n32_adj_388)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i17_4_lut_adj_564 (.A(addr[13]), .B(addr[6]), .C(addr[11]), .D(addr[15]), 
         .Z(n46_adj_389)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut_adj_564.init = 16'hfffe;
    LUT4 i15_3_lut (.A(addr[22]), .B(addr[21]), .C(addr[10]), .Z(n44_adj_390)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15_3_lut.init = 16'hfefe;
    LUT4 i23_4_lut (.A(addr[7]), .B(n46_adj_389), .C(n32_adj_388), .D(addr[17]), 
         .Z(n52_adj_391)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i25_4_lut (.A(addr[3]), .B(n50_adj_386), .C(n40_adj_385), .D(addr[4]), 
         .Z(n54_adj_392)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i25_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut_adj_565 (.A(addr[16]), .B(n48), .C(n36_adj_387), .D(addr[18]), 
         .Z(n53)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut_adj_565.init = 16'hfffe;
    LUT4 i26_4_lut_adj_566 (.A(addr[26]), .B(n52_adj_391), .C(n44_adj_390), 
         .D(addr[30]), .Z(n55_adj_393)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26_4_lut_adj_566.init = 16'hfffe;
    LUT4 i1_4_lut_adj_567 (.A(n55_adj_393), .B(addr[31]), .C(n53), .D(n54_adj_392), 
         .Z(n65)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_567.init = 16'hcccd;
    CCU2D equal_232_0 (.A0(n[31]), .B0(n3921), .C0(GND_net), .D0(GND_net), 
          .A1(n[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n60985));
    defparam equal_232_0.INIT0 = 16'h9000;
    defparam equal_232_0.INIT1 = 16'haaaa;
    defparam equal_232_0.INJECT1_0 = "NO";
    defparam equal_232_0.INJECT1_1 = "YES";
    CCU2D equal_152_32 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n60984), 
          .S0(n2664));
    defparam equal_152_32.INIT0 = 16'hFFFF;
    defparam equal_152_32.INIT1 = 16'h0000;
    defparam equal_152_32.INJECT1_0 = "NO";
    defparam equal_152_32.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_33 (.A0(i_c[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62189), 
          .S0(n134_adj_409[31]));
    defparam i_4655_add_4_33.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_33.INIT1 = 16'h0000;
    defparam i_4655_add_4_33.INJECT1_0 = "NO";
    defparam i_4655_add_4_33.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_31 (.A0(i_c[29]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62188), 
          .COUT(n62189), .S0(n134_adj_409[29]), .S1(n134_adj_409[30]));
    defparam i_4655_add_4_31.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_31.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_31.INJECT1_0 = "NO";
    defparam i_4655_add_4_31.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_29 (.A0(i_c[27]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62187), 
          .COUT(n62188), .S0(n134_adj_409[27]), .S1(n134_adj_409[28]));
    defparam i_4655_add_4_29.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_29.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_29.INJECT1_0 = "NO";
    defparam i_4655_add_4_29.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_27 (.A0(i_c[25]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62186), 
          .COUT(n62187), .S0(n134_adj_409[25]), .S1(n134_adj_409[26]));
    defparam i_4655_add_4_27.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_27.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_27.INJECT1_0 = "NO";
    defparam i_4655_add_4_27.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_25 (.A0(i_c[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62185), 
          .COUT(n62186), .S0(n134_adj_409[23]), .S1(n134_adj_409[24]));
    defparam i_4655_add_4_25.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_25.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_25.INJECT1_0 = "NO";
    defparam i_4655_add_4_25.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_23 (.A0(i_c[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62184), 
          .COUT(n62185), .S0(n134_adj_409[21]), .S1(n134_adj_409[22]));
    defparam i_4655_add_4_23.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_23.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_23.INJECT1_0 = "NO";
    defparam i_4655_add_4_23.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_21 (.A0(i_c[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62183), 
          .COUT(n62184), .S0(n134_adj_409[19]), .S1(n134_adj_409[20]));
    defparam i_4655_add_4_21.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_21.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_21.INJECT1_0 = "NO";
    defparam i_4655_add_4_21.INJECT1_1 = "NO";
    LUT4 mux_141_Mux_1_i7_4_lut (.A(n67359), .B(\hidden_outputs[4] [1]), 
         .C(h[2]), .D(n70861), .Z(n2448[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_1_i7_4_lut.init = 16'h0aca;
    CCU2D i_4655_add_4_19 (.A0(i_c[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62182), 
          .COUT(n62183), .S0(n134_adj_409[17]), .S1(n134_adj_409[18]));
    defparam i_4655_add_4_19.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_19.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_19.INJECT1_0 = "NO";
    defparam i_4655_add_4_19.INJECT1_1 = "NO";
    LUT4 mux_237_Mux_1_i1_3_lut (.A(\mlp_outputs[0] [1]), .B(\mlp_outputs[1] [1]), 
         .C(o[0]), .Z(n4478[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_1_i1_3_lut.init = 16'hcaca;
    CCU2D i_4655_add_4_17 (.A0(i_c[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62181), 
          .COUT(n62182), .S0(n134_adj_409[15]), .S1(n134_adj_409[16]));
    defparam i_4655_add_4_17.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_17.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_17.INJECT1_0 = "NO";
    defparam i_4655_add_4_17.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_15 (.A0(i_c[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i_c[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62180), 
          .COUT(n62181), .S0(n134_adj_409[13]), .S1(n134_adj_409[14]));
    defparam i_4655_add_4_15.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_15.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_15.INJECT1_0 = "NO";
    defparam i_4655_add_4_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_568 (.A(n2448[1]), .B(n23104), .Z(n22793)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_568.init = 16'h8888;
    LUT4 i2_4_lut_adj_569 (.A(n22793), .B(n22796), .C(weight[1]), .D(n70860), 
         .Z(n62966)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_569.init = 16'hfeee;
    CCU2D i_4655_add_4_13 (.A0(\i[11] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\i[12] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62179), 
          .COUT(n62180), .S0(n134_adj_409[11]), .S1(n134_adj_409[12]));
    defparam i_4655_add_4_13.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_13.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_13.INJECT1_0 = "NO";
    defparam i_4655_add_4_13.INJECT1_1 = "NO";
    LUT4 mux_141_Mux_2_i7_4_lut (.A(n67362), .B(\hidden_outputs[4] [2]), 
         .C(h[2]), .D(n70861), .Z(n2448[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_2_i7_4_lut.init = 16'h0aca;
    CCU2D i_4655_add_4_11 (.A0(\i[9] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62178), 
          .COUT(n62179), .S0(n134_adj_409[9]), .S1(n134_adj_409[10]));
    defparam i_4655_add_4_11.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_11.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_11.INJECT1_0 = "NO";
    defparam i_4655_add_4_11.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_9 (.A0(\i[7] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\i[8] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62177), 
          .COUT(n62178), .S0(n134_adj_409[7]), .S1(n134_adj_409[8]));
    defparam i_4655_add_4_9.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_9.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_9.INJECT1_0 = "NO";
    defparam i_4655_add_4_9.INJECT1_1 = "NO";
    LUT4 mux_237_Mux_2_i1_3_lut (.A(\mlp_outputs[0] [2]), .B(\mlp_outputs[1] [2]), 
         .C(o[0]), .Z(n4478[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_2_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_570 (.A(n2448[2]), .B(n23104), .Z(n22784)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_570.init = 16'h8888;
    LUT4 i2_4_lut_adj_571 (.A(n22784), .B(n22787), .C(weight[2]), .D(n70860), 
         .Z(n62964)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_571.init = 16'hfeee;
    LUT4 mux_141_Mux_3_i7_4_lut (.A(n67365), .B(\hidden_outputs[4] [3]), 
         .C(h[2]), .D(n70861), .Z(n2448[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_3_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_3_i1_3_lut (.A(\mlp_outputs[0] [3]), .B(\mlp_outputs[1] [3]), 
         .C(o[0]), .Z(n4478[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_572 (.A(n2448[3]), .B(n23104), .Z(n23123)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_572.init = 16'h8888;
    LUT4 i2_4_lut_adj_573 (.A(n23123), .B(n23126), .C(weight[3]), .D(n70860), 
         .Z(n63150)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_573.init = 16'hfeee;
    LUT4 mux_141_Mux_4_i7_4_lut (.A(n67368), .B(\hidden_outputs[4] [4]), 
         .C(h[2]), .D(n70861), .Z(n2448[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_4_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_4_i1_3_lut (.A(\mlp_outputs[0] [4]), .B(\mlp_outputs[1] [4]), 
         .C(o[0]), .Z(n4478[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_574 (.A(n2448[4]), .B(n23104), .Z(n23114)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_574.init = 16'h8888;
    LUT4 i2_4_lut_adj_575 (.A(n23114), .B(n23117), .C(weight[4]), .D(n70860), 
         .Z(n63147)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_575.init = 16'hfeee;
    LUT4 mux_141_Mux_5_i7_4_lut (.A(n67371), .B(\hidden_outputs[4] [5]), 
         .C(h[2]), .D(n70861), .Z(n2448[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_5_i7_4_lut.init = 16'h0aca;
    CCU2D i_4655_add_4_7 (.A0(\i[5] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\i[6] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62176), 
          .COUT(n62177), .S0(n134_adj_409[5]), .S1(n134_adj_409[6]));
    defparam i_4655_add_4_7.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_7.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_7.INJECT1_0 = "NO";
    defparam i_4655_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_237_Mux_5_i1_3_lut (.A(\mlp_outputs[0] [5]), .B(\mlp_outputs[1] [5]), 
         .C(o[0]), .Z(n4478[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_5_i1_3_lut.init = 16'hcaca;
    CCU2D i_4655_add_4_5 (.A0(\i[3] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\i[4] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62175), 
          .COUT(n62176), .S0(n134_adj_409[3]), .S1(n134_adj_409[4]));
    defparam i_4655_add_4_5.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_5.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_5.INJECT1_0 = "NO";
    defparam i_4655_add_4_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_576 (.A(n2448[5]), .B(n23104), .Z(n23105)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_576.init = 16'h8888;
    LUT4 i2_4_lut_adj_577 (.A(n23105), .B(n23108), .C(weight[5]), .D(n70860), 
         .Z(n63139)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_577.init = 16'hfeee;
    LUT4 mux_141_Mux_6_i7_4_lut (.A(n67374), .B(\hidden_outputs[4] [6]), 
         .C(h[2]), .D(n70861), .Z(n2448[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_6_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_6_i1_3_lut (.A(\mlp_outputs[0] [6]), .B(\mlp_outputs[1] [6]), 
         .C(o[0]), .Z(n4478[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_6_i1_3_lut.init = 16'hcaca;
    CCU2D i_4655_add_4_3 (.A0(i[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62174), 
          .COUT(n62175), .S0(n134_adj_409[1]), .S1(n134_adj_409[2]));
    defparam i_4655_add_4_3.INIT0 = 16'hfaaa;
    defparam i_4655_add_4_3.INIT1 = 16'hfaaa;
    defparam i_4655_add_4_3.INJECT1_0 = "NO";
    defparam i_4655_add_4_3.INJECT1_1 = "NO";
    CCU2D i_4655_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(i[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62174), 
          .S1(n134_adj_409[0]));
    defparam i_4655_add_4_1.INIT0 = 16'hF000;
    defparam i_4655_add_4_1.INIT1 = 16'h0555;
    defparam i_4655_add_4_1.INJECT1_0 = "NO";
    defparam i_4655_add_4_1.INJECT1_1 = "NO";
    CCU2D equal_152_32_49660 (.A0(h[7]), .B0(h[6]), .C0(h[5]), .D0(h[4]), 
          .A1(h[4]), .B1(h[3]), .C1(h[2]), .D1(h[1]), .CIN(n60983), 
          .COUT(n60984));
    defparam equal_152_32_49660.INIT0 = 16'h8001;
    defparam equal_152_32_49660.INIT1 = 16'h8001;
    defparam equal_152_32_49660.INJECT1_0 = "YES";
    defparam equal_152_32_49660.INJECT1_1 = "YES";
    LUT4 i1_2_lut_adj_578 (.A(n2448[6]), .B(n23104), .Z(n23096)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_578.init = 16'h8888;
    LUT4 i2_4_lut_adj_579 (.A(n23096), .B(n23099), .C(weight[6]), .D(n70860), 
         .Z(n63131)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_579.init = 16'hfeee;
    LUT4 mux_141_Mux_7_i7_4_lut (.A(n67377), .B(\hidden_outputs[4] [7]), 
         .C(h[2]), .D(n70861), .Z(n2448[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_7_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_7_i1_3_lut (.A(\mlp_outputs[0] [7]), .B(\mlp_outputs[1] [7]), 
         .C(o[0]), .Z(n4478[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_580 (.A(n2448[7]), .B(n23104), .Z(n23087)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_580.init = 16'h8888;
    LUT4 i2_4_lut_adj_581 (.A(n23087), .B(n23090), .C(weight[7]), .D(n70860), 
         .Z(n63128)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_581.init = 16'hfeee;
    LUT4 mux_141_Mux_8_i7_4_lut (.A(n67380), .B(\hidden_outputs[4] [8]), 
         .C(h[2]), .D(n70861), .Z(n2448[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_8_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_8_i1_3_lut (.A(\mlp_outputs[0] [8]), .B(\mlp_outputs[1] [8]), 
         .C(o[0]), .Z(n4478[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_8_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_582 (.A(n2448[8]), .B(n23104), .Z(n23078)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_582.init = 16'h8888;
    LUT4 i2_4_lut_adj_583 (.A(n23078), .B(n23081), .C(weight[8]), .D(n70860), 
         .Z(n63122)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_583.init = 16'hfeee;
    LUT4 mux_141_Mux_9_i7_4_lut (.A(n67383), .B(\hidden_outputs[4] [9]), 
         .C(h[2]), .D(n70861), .Z(n2448[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_9_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_9_i1_3_lut (.A(\mlp_outputs[0] [9]), .B(\mlp_outputs[1] [9]), 
         .C(o[0]), .Z(n4478[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_9_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_584 (.A(n2448[9]), .B(n23104), .Z(n23069)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_584.init = 16'h8888;
    LUT4 i2_4_lut_adj_585 (.A(n23069), .B(n23072), .C(weight[9]), .D(n70860), 
         .Z(n63120)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_585.init = 16'hfeee;
    LUT4 mux_141_Mux_10_i7_4_lut (.A(n67386), .B(\hidden_outputs[4] [10]), 
         .C(h[2]), .D(n70861), .Z(n2448[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_10_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_10_i1_3_lut (.A(\mlp_outputs[0] [10]), .B(\mlp_outputs[1] [10]), 
         .C(o[0]), .Z(n4478[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_10_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_586 (.A(n2448[10]), .B(n23104), .Z(n23060)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_586.init = 16'h8888;
    LUT4 i2_4_lut_adj_587 (.A(n23060), .B(n23063), .C(weight[10]), .D(n70860), 
         .Z(n63116)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_587.init = 16'hfeee;
    LUT4 mux_141_Mux_11_i7_4_lut (.A(n67389), .B(\hidden_outputs[4] [11]), 
         .C(h[2]), .D(n70861), .Z(n2448[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_11_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_11_i1_3_lut (.A(\mlp_outputs[0] [11]), .B(\mlp_outputs[1] [11]), 
         .C(o[0]), .Z(n4478[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_11_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_588 (.A(n2448[11]), .B(n23104), .Z(n23051)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_588.init = 16'h8888;
    LUT4 i2_4_lut_adj_589 (.A(n23051), .B(n23054), .C(weight[11]), .D(n70860), 
         .Z(n63115)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_589.init = 16'hfeee;
    LUT4 mux_141_Mux_12_i7_4_lut (.A(n67392), .B(\hidden_outputs[4] [12]), 
         .C(h[2]), .D(n70861), .Z(n2448[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_12_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_12_i1_3_lut (.A(\mlp_outputs[0] [12]), .B(\mlp_outputs[1] [12]), 
         .C(o[0]), .Z(n4478[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_12_i1_3_lut.init = 16'hcaca;
    CCU2D equal_152_30 (.A0(h[13]), .B0(h[12]), .C0(h[11]), .D0(h[10]), 
          .A1(h[10]), .B1(h[9]), .C1(h[8]), .D1(h[7]), .CIN(n60982), 
          .COUT(n60983));
    defparam equal_152_30.INIT0 = 16'h8001;
    defparam equal_152_30.INIT1 = 16'h8001;
    defparam equal_152_30.INJECT1_0 = "YES";
    defparam equal_152_30.INJECT1_1 = "YES";
    LUT4 i1_2_lut_adj_590 (.A(n2448[12]), .B(n23104), .Z(n23033)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_590.init = 16'h8888;
    LUT4 i2_4_lut_adj_591 (.A(n23033), .B(n23036), .C(weight[12]), .D(n70860), 
         .Z(n63109)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_591.init = 16'hfeee;
    LUT4 mux_141_Mux_13_i7_4_lut (.A(n67395), .B(\hidden_outputs[4] [13]), 
         .C(h[2]), .D(n70861), .Z(n2448[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_13_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_13_i1_3_lut (.A(\mlp_outputs[0] [13]), .B(\mlp_outputs[1] [13]), 
         .C(o[0]), .Z(n4478[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_13_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_592 (.A(n2448[13]), .B(n23104), .Z(n23042)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_592.init = 16'h8888;
    LUT4 i2_4_lut_adj_593 (.A(n23042), .B(n23045), .C(weight[13]), .D(n70860), 
         .Z(n63114)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_593.init = 16'hfeee;
    LUT4 mux_141_Mux_14_i7_4_lut (.A(n67398), .B(\hidden_outputs[4] [14]), 
         .C(h[2]), .D(n70861), .Z(n2448[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_14_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_14_i1_3_lut (.A(\mlp_outputs[0] [14]), .B(\mlp_outputs[1] [14]), 
         .C(o[0]), .Z(n4478[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_14_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_594 (.A(n2448[14]), .B(n23104), .Z(n23024)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_594.init = 16'h8888;
    LUT4 i2_4_lut_adj_595 (.A(n23024), .B(n23027), .C(weight[14]), .D(n70860), 
         .Z(n63107)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_595.init = 16'hfeee;
    LUT4 mux_141_Mux_15_i7_4_lut (.A(n67401), .B(\hidden_outputs[4] [15]), 
         .C(h[2]), .D(n70861), .Z(n2448[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_15_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_15_i1_3_lut (.A(\mlp_outputs[0] [15]), .B(\mlp_outputs[1] [15]), 
         .C(o[0]), .Z(n4478[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_15_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_596 (.A(n2448[15]), .B(n23104), .Z(n23006)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_596.init = 16'h8888;
    LUT4 i2_4_lut_adj_597 (.A(n23006), .B(n23009), .C(weight[15]), .D(n70860), 
         .Z(n63105)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_597.init = 16'hfeee;
    LUT4 mux_141_Mux_16_i7_4_lut (.A(n67404), .B(\hidden_outputs[4] [16]), 
         .C(h[2]), .D(n70861), .Z(n2448[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_16_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_16_i1_3_lut (.A(\mlp_outputs[0] [16]), .B(\mlp_outputs[1] [16]), 
         .C(o[0]), .Z(n4478[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_16_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_598 (.A(n2448[16]), .B(n23104), .Z(n23015)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_598.init = 16'h8888;
    LUT4 i2_4_lut_adj_599 (.A(n23015), .B(n23018), .C(weight[16]), .D(n70860), 
         .Z(n63106)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_599.init = 16'hfeee;
    LUT4 mux_141_Mux_17_i7_4_lut (.A(n67407), .B(\hidden_outputs[4] [17]), 
         .C(h[2]), .D(n70861), .Z(n2448[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_17_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_17_i1_3_lut (.A(\mlp_outputs[0] [17]), .B(\mlp_outputs[1] [17]), 
         .C(o[0]), .Z(n4478[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_17_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_600 (.A(n2448[17]), .B(n23104), .Z(n22997)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_600.init = 16'h8888;
    LUT4 i2_4_lut_adj_601 (.A(n22997), .B(n23000), .C(weight[17]), .D(n70860), 
         .Z(n63104)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_601.init = 16'hfeee;
    LUT4 mux_141_Mux_18_i7_4_lut (.A(n67410), .B(\hidden_outputs[4] [18]), 
         .C(h[2]), .D(n70861), .Z(n2448[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_18_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_18_i1_3_lut (.A(\mlp_outputs[0] [18]), .B(\mlp_outputs[1] [18]), 
         .C(o[0]), .Z(n4478[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_18_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_602 (.A(n2448[18]), .B(n23104), .Z(n22988)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_602.init = 16'h8888;
    LUT4 i2_4_lut_adj_603 (.A(n22988), .B(n22991), .C(weight[18]), .D(n70860), 
         .Z(n63103)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_603.init = 16'hfeee;
    LUT4 mux_141_Mux_19_i7_4_lut (.A(n67413), .B(\hidden_outputs[4] [19]), 
         .C(h[2]), .D(n70861), .Z(n2448[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_19_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_19_i1_3_lut (.A(\mlp_outputs[0] [19]), .B(\mlp_outputs[1] [19]), 
         .C(o[0]), .Z(n4478[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_19_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_604 (.A(n2448[19]), .B(n23104), .Z(n22979)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_604.init = 16'h8888;
    LUT4 i2_4_lut_adj_605 (.A(n22979), .B(n22982), .C(weight[19]), .D(n70860), 
         .Z(n63102)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_605.init = 16'hfeee;
    LUT4 mux_141_Mux_20_i7_4_lut (.A(n67416), .B(\hidden_outputs[4] [20]), 
         .C(h[2]), .D(n70861), .Z(n2448[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_20_i7_4_lut.init = 16'h0aca;
    CCU2D equal_152_28 (.A0(h[19]), .B0(h[18]), .C0(h[17]), .D0(h[16]), 
          .A1(h[16]), .B1(h[15]), .C1(h[14]), .D1(h[13]), .CIN(n60981), 
          .COUT(n60982));
    defparam equal_152_28.INIT0 = 16'h8001;
    defparam equal_152_28.INIT1 = 16'h8001;
    defparam equal_152_28.INJECT1_0 = "YES";
    defparam equal_152_28.INJECT1_1 = "YES";
    LUT4 mux_237_Mux_20_i1_3_lut (.A(\mlp_outputs[0] [20]), .B(\mlp_outputs[1] [20]), 
         .C(o[0]), .Z(n4478[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_20_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_606 (.A(n2448[20]), .B(n23104), .Z(n22766)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_606.init = 16'h8888;
    LUT4 i2_4_lut_adj_607 (.A(n22766), .B(n22769), .C(weight[20]), .D(n70860), 
         .Z(n62961)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_607.init = 16'hfeee;
    LUT4 mux_141_Mux_21_i7_4_lut (.A(n67419), .B(\hidden_outputs[4] [21]), 
         .C(h[2]), .D(n70861), .Z(n2448[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_21_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_21_i1_3_lut (.A(\mlp_outputs[0] [21]), .B(\mlp_outputs[1] [21]), 
         .C(o[0]), .Z(n4478[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_21_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_608 (.A(n2448[21]), .B(n23104), .Z(n22970)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_608.init = 16'h8888;
    LUT4 i2_4_lut_adj_609 (.A(n22970), .B(n22973), .C(weight[21]), .D(n70860), 
         .Z(n63070)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_609.init = 16'hfeee;
    LUT4 mux_141_Mux_22_i7_4_lut (.A(n67422), .B(\hidden_outputs[4] [22]), 
         .C(h[2]), .D(n70861), .Z(n2448[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_22_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_22_i1_3_lut (.A(\mlp_outputs[0] [22]), .B(\mlp_outputs[1] [22]), 
         .C(o[0]), .Z(n4478[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_22_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_610 (.A(n2448[22]), .B(n23104), .Z(n22961)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_610.init = 16'h8888;
    LUT4 i2_4_lut_adj_611 (.A(n22961), .B(n22964), .C(weight[22]), .D(n70860), 
         .Z(n63069)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_611.init = 16'hfeee;
    LUT4 mux_237_Mux_23_i1_3_lut (.A(\mlp_outputs[0] [23]), .B(\mlp_outputs[1] [23]), 
         .C(o[0]), .Z(n4478[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_23_i1_3_lut.init = 16'hcaca;
    LUT4 mux_141_Mux_23_i7_4_lut (.A(n67425), .B(\hidden_outputs[4] [23]), 
         .C(h[2]), .D(n70861), .Z(n2448[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_23_i7_4_lut.init = 16'h0aca;
    LUT4 i2_4_lut_adj_612 (.A(n2448[23]), .B(n4478[23]), .C(n23104), .D(n70813), 
         .Z(n6_adj_394)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_612.init = 16'heca0;
    LUT4 i3_4_lut_adj_613 (.A(weight[23]), .B(n6_adj_394), .C(n22276), 
         .D(n70860), .Z(n63156)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut_adj_613.init = 16'hfefc;
    LUT4 mux_237_Mux_25_i1_3_lut (.A(\mlp_outputs[0] [25]), .B(\mlp_outputs[1] [25]), 
         .C(o[0]), .Z(n4478[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_25_i1_3_lut.init = 16'hcaca;
    LUT4 mux_141_Mux_25_i7_4_lut (.A(n67431), .B(\hidden_outputs[4] [25]), 
         .C(h[2]), .D(n70861), .Z(n2448[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_25_i7_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_614 (.A(weight[25]), .B(n2448[25]), .C(n70860), 
         .D(n23104), .Z(n4_adj_395)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_614.init = 16'heca0;
    LUT4 i1_4_lut_adj_615 (.A(n22276), .B(n4478[25]), .C(n4_adj_395), 
         .D(n70813), .Z(n66524)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_615.init = 16'hfefa;
    LUT4 mux_237_Mux_27_i1_3_lut (.A(\mlp_outputs[0] [27]), .B(\mlp_outputs[1] [27]), 
         .C(o[0]), .Z(n4478[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_27_i1_3_lut.init = 16'hcaca;
    LUT4 mux_141_Mux_27_i7_4_lut (.A(n67437), .B(\hidden_outputs[4] [27]), 
         .C(h[2]), .D(n70861), .Z(n2448[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_27_i7_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_616 (.A(weight[27]), .B(n2448[27]), .C(n70860), 
         .D(n23104), .Z(n4_adj_396)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_616.init = 16'heca0;
    LUT4 i1_4_lut_adj_617 (.A(n22276), .B(n4478[27]), .C(n4_adj_396), 
         .D(n70813), .Z(n66522)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_617.init = 16'hfefa;
    LUT4 mux_141_Mux_30_i7_4_lut (.A(n67446), .B(\hidden_outputs[4] [30]), 
         .C(h[2]), .D(n70861), .Z(n2448[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_30_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_30_i1_3_lut (.A(\mlp_outputs[0] [30]), .B(\mlp_outputs[1] [30]), 
         .C(o[0]), .Z(n4478[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_30_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_618 (.A(n2448[30]), .B(n23104), .Z(n22754)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_618.init = 16'h8888;
    LUT4 i2_4_lut_adj_619 (.A(n22754), .B(n22757), .C(weight[30]), .D(n70860), 
         .Z(n62958)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_619.init = 16'hfeee;
    LUT4 mux_141_Mux_31_i7_4_lut (.A(n67449), .B(\hidden_outputs[4] [31]), 
         .C(h[2]), .D(n70861), .Z(n2448[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam mux_141_Mux_31_i7_4_lut.init = 16'h0aca;
    LUT4 mux_237_Mux_31_i1_3_lut (.A(\mlp_outputs[0] [31]), .B(\mlp_outputs[1] [31]), 
         .C(o[0]), .Z(n3998[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_237_Mux_31_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_620 (.A(n2448[31]), .B(n23104), .Z(n22952)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_620.init = 16'h8888;
    LUT4 i2_4_lut_adj_621 (.A(n22952), .B(n22955), .C(weight[31]), .D(n70860), 
         .Z(n63068)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_621.init = 16'hfeee;
    CCU2D equal_152_26 (.A0(h[25]), .B0(h[24]), .C0(h[23]), .D0(h[22]), 
          .A1(h[22]), .B1(h[21]), .C1(h[20]), .D1(h[19]), .CIN(n60980), 
          .COUT(n60981));
    defparam equal_152_26.INIT0 = 16'h8001;
    defparam equal_152_26.INIT1 = 16'h8001;
    defparam equal_152_26.INJECT1_0 = "YES";
    defparam equal_152_26.INJECT1_1 = "YES";
    LUT4 i54378_3_lut (.A(\temp_outputs[2] [24]), .B(\temp_outputs[3] [24]), 
         .C(i[0]), .Z(n67289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54378_3_lut.init = 16'hcaca;
    LUT4 i54377_3_lut (.A(\temp_outputs[0] [24]), .B(\temp_outputs[1] [24]), 
         .C(i[0]), .Z(n67288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54377_3_lut.init = 16'hcaca;
    LUT4 i10011_1_lut_2_lut (.A(n14054), .B(numL[0]), .Z(n3921)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i10011_1_lut_2_lut.init = 16'h9999;
    LUT4 i1_2_lut_rep_897 (.A(n14054), .B(numL[0]), .Z(n70867)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_897.init = 16'h6666;
    LUT4 i1_4_lut_adj_622 (.A(n11102[10]), .B(n61278[10]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_397)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_622.init = 16'heca0;
    LUT4 i2_4_lut_adj_623 (.A(n61250[10]), .B(addr[10]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_398)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_623.init = 16'heca0;
    LUT4 i4_4_lut_adj_624 (.A(n7_adj_398), .B(n61312[10]), .C(n6_adj_397), 
         .D(n2022[32]), .Z(n63119)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_624.init = 16'hfefa;
    LUT4 i54375_3_lut (.A(\temp_outputs[2] [25]), .B(\temp_outputs[3] [25]), 
         .C(i[0]), .Z(n67286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54375_3_lut.init = 16'hcaca;
    LUT4 i54374_3_lut (.A(\temp_outputs[0] [25]), .B(\temp_outputs[1] [25]), 
         .C(i[0]), .Z(n67285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54374_3_lut.init = 16'hcaca;
    LUT4 i54372_3_lut (.A(\temp_outputs[2] [26]), .B(\temp_outputs[3] [26]), 
         .C(i[0]), .Z(n67283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54372_3_lut.init = 16'hcaca;
    LUT4 i54371_3_lut (.A(\temp_outputs[0] [26]), .B(\temp_outputs[1] [26]), 
         .C(i[0]), .Z(n67282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54371_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_625 (.A(n11102[11]), .B(n61278[11]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_399)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_625.init = 16'heca0;
    LUT4 i2_4_lut_adj_626 (.A(n61250[11]), .B(addr[11]), .C(n2022[10]), 
         .D(n2022[1]), .Z(n7_adj_400)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_626.init = 16'heca0;
    LUT4 i4_4_lut_adj_627 (.A(n7_adj_400), .B(n61312[11]), .C(n6_adj_399), 
         .D(n2022[32]), .Z(n63155)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i4_4_lut_adj_627.init = 16'hfefa;
    LUT4 i1_4_lut_adj_628 (.A(\mlp_outputs[0] [1]), .B(n70809), .C(float_alu_c[1]), 
         .D(o[0]), .Z(n23426)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_628.init = 16'h88c0;
    LUT4 i2_4_lut_adj_629 (.A(n23426), .B(n32_adj_73), .C(\mlp_outputs[0] [1]), 
         .D(n2022[39]), .Z(n63213)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_629.init = 16'hfeee;
    LUT4 i1_4_lut_adj_630 (.A(\mlp_outputs[0] [2]), .B(n70809), .C(float_alu_c[2]), 
         .D(o[0]), .Z(n23402)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_630.init = 16'h88c0;
    LUT4 i2_4_lut_adj_631 (.A(n23402), .B(n32_adj_74), .C(\mlp_outputs[0] [2]), 
         .D(n2022[39]), .Z(n63203)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_631.init = 16'hfeee;
    LUT4 i1_4_lut_adj_632 (.A(\mlp_outputs[0] [3]), .B(n70809), .C(float_alu_c[3]), 
         .D(o[0]), .Z(n23408)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_632.init = 16'h88c0;
    LUT4 i2_4_lut_adj_633 (.A(n23408), .B(n32_adj_75), .C(\mlp_outputs[0] [3]), 
         .D(n2022[39]), .Z(n63206)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_633.init = 16'hfeee;
    LUT4 i1_4_lut_adj_634 (.A(\mlp_outputs[0] [4]), .B(n70809), .C(float_alu_c[4]), 
         .D(o[0]), .Z(n22877)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_634.init = 16'h88c0;
    LUT4 i2_4_lut_adj_635 (.A(n32_adj_76), .B(n22877), .C(\mlp_outputs[0] [4]), 
         .D(n2022[39]), .Z(n62990)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_635.init = 16'hfeee;
    LUT4 i1_4_lut_adj_636 (.A(\mlp_outputs[0] [5]), .B(n70809), .C(float_alu_c[5]), 
         .D(o[0]), .Z(n23423)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_636.init = 16'h88c0;
    LUT4 i1_4_lut_adj_637 (.A(n32_adj_80), .B(\mlp_outputs[0] [5]), .C(n23423), 
         .D(n2022[39]), .Z(n66368)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_637.init = 16'hfefa;
    LUT4 i1_4_lut_adj_638 (.A(\mlp_outputs[0] [6]), .B(n70809), .C(float_alu_c[6]), 
         .D(o[0]), .Z(n23480)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_638.init = 16'h88c0;
    LUT4 i1_4_lut_adj_639 (.A(n32_adj_84), .B(\mlp_outputs[0] [6]), .C(n23480), 
         .D(n2022[39]), .Z(n66350)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_639.init = 16'hfefa;
    LUT4 i1_4_lut_adj_640 (.A(\mlp_outputs[0] [7]), .B(n70809), .C(float_alu_c[7]), 
         .D(o[0]), .Z(n22817)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_640.init = 16'h88c0;
    LUT4 i2_4_lut_adj_641 (.A(n32_adj_91), .B(n22817), .C(\mlp_outputs[0] [7]), 
         .D(n2022[39]), .Z(n62972)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_641.init = 16'hfeee;
    LUT4 i1_4_lut_adj_642 (.A(\mlp_outputs[0] [8]), .B(n70809), .C(float_alu_c[8]), 
         .D(o[0]), .Z(n23486)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_642.init = 16'h88c0;
    LUT4 i2_4_lut_adj_643 (.A(n23486), .B(n32_adj_92), .C(\mlp_outputs[0] [8]), 
         .D(n2022[39]), .Z(n63235)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_643.init = 16'hfeee;
    LUT4 i1_4_lut_adj_644 (.A(\mlp_outputs[0] [9]), .B(n70809), .C(float_alu_c[9]), 
         .D(o[0]), .Z(n22823)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_644.init = 16'h88c0;
    LUT4 i1_4_lut_adj_645 (.A(n32_adj_93), .B(n22823), .C(\mlp_outputs[0] [9]), 
         .D(n2022[39]), .Z(n66446)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_645.init = 16'hfeee;
    LUT4 i1_4_lut_adj_646 (.A(\mlp_outputs[0] [10]), .B(n70809), .C(float_alu_c[10]), 
         .D(o[0]), .Z(n23471)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_646.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_647 (.A(n2022[24]), .B(n2022[22]), .C(n2448[26]), 
         .Z(n22925)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_647.init = 16'he0e0;
    LUT4 i1_2_lut_3_lut_adj_648 (.A(n2022[24]), .B(n2022[22]), .C(n2448[25]), 
         .Z(n22922)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_648.init = 16'he0e0;
    LUT4 i1_4_lut_adj_649 (.A(n32_adj_94), .B(\mlp_outputs[0] [10]), .C(n23471), 
         .D(n2022[39]), .Z(n66342)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_649.init = 16'hfefa;
    LUT4 i1_2_lut_3_lut_adj_650 (.A(n2022[24]), .B(n2022[22]), .C(n2448[23]), 
         .Z(n22919)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_650.init = 16'he0e0;
    LUT4 i1_4_lut_adj_651 (.A(\mlp_outputs[0] [11]), .B(n70809), .C(float_alu_c[11]), 
         .D(o[0]), .Z(n22586)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_651.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_652 (.A(n2022[24]), .B(n2022[22]), .C(n2448[27]), 
         .Z(n22934)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_652.init = 16'he0e0;
    LUT4 i1_4_lut_adj_653 (.A(n32_adj_95), .B(n22586), .C(\mlp_outputs[0] [11]), 
         .D(n2022[39]), .Z(n66396)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_653.init = 16'hfeee;
    LUT4 i1_4_lut_adj_654 (.A(\mlp_outputs[0] [12]), .B(n70809), .C(float_alu_c[12]), 
         .D(o[0]), .Z(n23477)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_654.init = 16'h88c0;
    LUT4 i2_4_lut_adj_655 (.A(n23477), .B(n32_adj_96), .C(\mlp_outputs[0] [12]), 
         .D(n2022[39]), .Z(n63232)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_655.init = 16'hfeee;
    LUT4 i1_4_lut_adj_656 (.A(\mlp_outputs[0] [13]), .B(n70809), .C(float_alu_c[13]), 
         .D(o[0]), .Z(n23468)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_656.init = 16'h88c0;
    LUT4 i2_4_lut_adj_657 (.A(n23468), .B(n32_adj_97), .C(\mlp_outputs[0] [13]), 
         .D(n2022[39]), .Z(n63227)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_657.init = 16'hfeee;
    CCU2D equal_152_24 (.A0(h[31]), .B0(h[30]), .C0(h[29]), .D0(h[28]), 
          .A1(h[28]), .B1(h[27]), .C1(h[26]), .D1(h[25]), .CIN(n60979), 
          .COUT(n60980));
    defparam equal_152_24.INIT0 = 16'h8001;
    defparam equal_152_24.INIT1 = 16'h8001;
    defparam equal_152_24.INJECT1_0 = "YES";
    defparam equal_152_24.INJECT1_1 = "YES";
    LUT4 i1_4_lut_adj_658 (.A(\mlp_outputs[0] [14]), .B(n70809), .C(float_alu_c[14]), 
         .D(o[0]), .Z(n22835)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_658.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_adj_659 (.A(n2022[24]), .B(n2022[22]), .C(n2448[29]), 
         .Z(n22931)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_659.init = 16'he0e0;
    LUT4 i1_4_lut_adj_660 (.A(n32_adj_98), .B(n22835), .C(\mlp_outputs[0] [14]), 
         .D(n2022[39]), .Z(n66442)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_660.init = 16'hfeee;
    LUT4 i3_2_lut_rep_894 (.A(n2022[24]), .B(n2022[22]), .Z(n70864)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_rep_894.init = 16'heeee;
    LUT4 i1_4_lut_adj_661 (.A(\mlp_outputs[0] [15]), .B(n70809), .C(float_alu_c[15]), 
         .D(o[0]), .Z(n23474)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_661.init = 16'h88c0;
    LUT4 i1_2_lut_rep_842_3_lut_4_lut (.A(n2022[37]), .B(n2022[46]), .C(n2022[35]), 
         .D(n2022[13]), .Z(n70812)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_842_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_662 (.A(n32_adj_99), .B(\mlp_outputs[0] [15]), .C(n23474), 
         .D(n2022[39]), .Z(n66320)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_662.init = 16'hfefa;
    LUT4 i1_2_lut_3_lut_4_lut_adj_663 (.A(n2022[37]), .B(n2022[46]), .C(n4478[28]), 
         .D(n70862), .Z(n23348)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_663.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_664 (.A(n2022[37]), .B(n2022[46]), .C(n4478[29]), 
         .D(n70862), .Z(n23528)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_664.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_665 (.A(n2022[37]), .B(n2022[46]), .C(n4478[0]), 
         .D(n70862), .Z(n22610)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_665.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_666 (.A(\mlp_outputs[0] [16]), .B(n70809), .C(float_alu_c[16]), 
         .D(o[0]), .Z(n22832)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_666.init = 16'h88c0;
    LUT4 i2_4_lut_adj_667 (.A(n32_adj_100), .B(n22832), .C(\mlp_outputs[0] [16]), 
         .D(n2022[39]), .Z(n62976)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_667.init = 16'hfeee;
    LUT4 i1_4_lut_adj_668 (.A(\mlp_outputs[0] [17]), .B(n70809), .C(float_alu_c[17]), 
         .D(o[0]), .Z(n23450)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_668.init = 16'h88c0;
    LUT4 i2_4_lut_adj_669 (.A(n23450), .B(n32_adj_101), .C(\mlp_outputs[0] [17]), 
         .D(n2022[39]), .Z(n63221)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_669.init = 16'hfeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_670 (.A(n2022[37]), .B(n2022[46]), .C(n3998[31]), 
         .D(n70862), .Z(n22955)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_670.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_671 (.A(\mlp_outputs[0] [18]), .B(n70809), .C(float_alu_c[18]), 
         .D(o[0]), .Z(n22838)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_671.init = 16'h88c0;
    LUT4 i2_4_lut_adj_672 (.A(n32_adj_102), .B(n22838), .C(\mlp_outputs[0] [18]), 
         .D(n2022[39]), .Z(n62978)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_672.init = 16'hfeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_673 (.A(n2022[37]), .B(n2022[46]), .C(n4478[30]), 
         .D(n70862), .Z(n22757)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_673.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_674 (.A(n2022[37]), .B(n2022[46]), .C(n4478[22]), 
         .D(n70862), .Z(n22964)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_674.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_675 (.A(\mlp_outputs[0] [19]), .B(n70809), .C(float_alu_c[19]), 
         .D(o[0]), .Z(n22844)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_675.init = 16'h88c0;
    LUT4 i1_4_lut_adj_676 (.A(n32_adj_103), .B(n22844), .C(\mlp_outputs[0] [19]), 
         .D(n2022[39]), .Z(n66440)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_676.init = 16'hfeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_677 (.A(n2022[37]), .B(n2022[46]), .C(n4478[21]), 
         .D(n70862), .Z(n22973)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_677.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_678 (.A(\mlp_outputs[0] [20]), .B(n70809), .C(float_alu_c[20]), 
         .D(o[0]), .Z(n23444)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_678.init = 16'h88c0;
    LUT4 i2_4_lut_adj_679 (.A(n23444), .B(n32_adj_105), .C(\mlp_outputs[0] [20]), 
         .D(n2022[39]), .Z(n63219)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_679.init = 16'hfeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_680 (.A(n2022[37]), .B(n2022[46]), .C(n4478[20]), 
         .D(n70862), .Z(n22769)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_680.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_681 (.A(\mlp_outputs[0] [21]), .B(n70809), .C(float_alu_c[21]), 
         .D(o[0]), .Z(n22847)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_681.init = 16'h88c0;
    LUT4 i1_4_lut_adj_682 (.A(n32_adj_106), .B(n22847), .C(\mlp_outputs[0] [21]), 
         .D(n2022[39]), .Z(n66438)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_682.init = 16'hfeee;
    LUT4 i1_4_lut_adj_683 (.A(\mlp_outputs[0] [22]), .B(n70809), .C(float_alu_c[22]), 
         .D(o[0]), .Z(n23441)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_683.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_684 (.A(n2022[37]), .B(n2022[46]), .C(n4478[19]), 
         .D(n70862), .Z(n22982)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_684.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_685 (.A(n2022[37]), .B(n2022[46]), .C(n4478[18]), 
         .D(n70862), .Z(n22991)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_685.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_686 (.A(n32_adj_107), .B(\mlp_outputs[0] [22]), .C(n23441), 
         .D(n2022[39]), .Z(n66362)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_686.init = 16'hfefa;
    LUT4 i1_2_lut_3_lut_4_lut_adj_687 (.A(n2022[37]), .B(n2022[46]), .C(n4478[17]), 
         .D(n70862), .Z(n23000)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_687.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_688 (.A(n2022[37]), .B(n2022[46]), .C(n4478[16]), 
         .D(n70862), .Z(n23018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_688.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_689 (.A(\mlp_outputs[0] [23]), .B(n70809), .C(float_alu_c[23]), 
         .D(o[0]), .Z(n22850)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_689.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_690 (.A(n2022[37]), .B(n2022[46]), .C(n4478[15]), 
         .D(n70862), .Z(n23009)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_690.init = 16'hf0e0;
    LUT4 i2_4_lut_adj_691 (.A(n32_adj_110), .B(n22850), .C(\mlp_outputs[0] [23]), 
         .D(n2022[39]), .Z(n62981)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_691.init = 16'hfeee;
    LUT4 i1_4_lut_adj_692 (.A(\mlp_outputs[0] [24]), .B(n70809), .C(float_alu_c[24]), 
         .D(o[0]), .Z(n23438)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_692.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_693 (.A(n2022[37]), .B(n2022[46]), .C(n4478[14]), 
         .D(n70862), .Z(n23027)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_693.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_694 (.A(n2022[37]), .B(n2022[46]), .C(n4478[13]), 
         .D(n70862), .Z(n23045)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_694.init = 16'hf0e0;
    LUT4 i2_4_lut_adj_695 (.A(n23438), .B(n32_adj_263), .C(\mlp_outputs[0] [24]), 
         .D(n2022[39]), .Z(n63217)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_695.init = 16'hfeee;
    LUT4 i1_4_lut_adj_696 (.A(\mlp_outputs[0] [25]), .B(n70809), .C(float_alu_c[25]), 
         .D(o[0]), .Z(n22853)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_696.init = 16'h88c0;
    LUT4 i1_4_lut_adj_697 (.A(n32_adj_270), .B(n22853), .C(\mlp_outputs[0] [25]), 
         .D(n2022[39]), .Z(n66436)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_697.init = 16'hfeee;
    LUT4 i1_4_lut_adj_698 (.A(\mlp_outputs[0] [26]), .B(n70809), .C(float_alu_c[26]), 
         .D(o[0]), .Z(n22856)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_698.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_699 (.A(n2022[37]), .B(n2022[46]), .C(n4478[12]), 
         .D(n70862), .Z(n23036)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_699.init = 16'hf0e0;
    LUT4 i2_4_lut_adj_700 (.A(n32_adj_280), .B(n22856), .C(\mlp_outputs[0] [26]), 
         .D(n2022[39]), .Z(n62983)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_700.init = 16'hfeee;
    LUT4 i1_4_lut_adj_701 (.A(\mlp_outputs[0] [27]), .B(n70809), .C(float_alu_c[27]), 
         .D(o[0]), .Z(n23432)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_701.init = 16'h88c0;
    LUT4 i2_4_lut_adj_702 (.A(n23432), .B(n32_adj_281), .C(\mlp_outputs[0] [27]), 
         .D(n2022[39]), .Z(n63215)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_702.init = 16'hfeee;
    LUT4 i1_4_lut_adj_703 (.A(\mlp_outputs[0] [28]), .B(n70809), .C(float_alu_c[28]), 
         .D(o[0]), .Z(n23429)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_703.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_704 (.A(n2022[37]), .B(n2022[46]), .C(n4478[11]), 
         .D(n70862), .Z(n23054)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_704.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_705 (.A(n32_adj_282), .B(\mlp_outputs[0] [28]), .C(n23429), 
         .D(n2022[39]), .Z(n66366)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_705.init = 16'hfefa;
    LUT4 i1_4_lut_adj_706 (.A(\mlp_outputs[0] [29]), .B(n70809), .C(float_alu_c[29]), 
         .D(o[0]), .Z(n22862)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_706.init = 16'h88c0;
    LUT4 i2_4_lut_adj_707 (.A(n32_adj_283), .B(n22862), .C(\mlp_outputs[0] [29]), 
         .D(n2022[39]), .Z(n62986)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_707.init = 16'hfeee;
    LUT4 i1_4_lut_adj_708 (.A(\mlp_outputs[0] [30]), .B(n70809), .C(float_alu_c[30]), 
         .D(o[0]), .Z(n23435)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_708.init = 16'h88c0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_709 (.A(n2022[37]), .B(n2022[46]), .C(n4478[10]), 
         .D(n70862), .Z(n23063)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_709.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_710 (.A(n2022[37]), .B(n2022[46]), .C(n4478[9]), 
         .D(n70862), .Z(n23072)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_710.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_711 (.A(n32_adj_285), .B(\mlp_outputs[0] [30]), .C(n23435), 
         .D(n2022[39]), .Z(n66364)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_711.init = 16'hfefa;
    LUT4 i54369_3_lut (.A(\temp_outputs[2] [27]), .B(\temp_outputs[3] [27]), 
         .C(i[0]), .Z(n67280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54369_3_lut.init = 16'hcaca;
    LUT4 i54368_3_lut (.A(\temp_outputs[0] [27]), .B(\temp_outputs[1] [27]), 
         .C(i[0]), .Z(n67279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54368_3_lut.init = 16'hcaca;
    CCU2D equal_152_0 (.A0(h[31]), .B0(n14054), .C0(GND_net), .D0(GND_net), 
          .A1(h[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n60979));
    defparam equal_152_0.INIT0 = 16'h9000;
    defparam equal_152_0.INIT1 = 16'haaaa;
    defparam equal_152_0.INJECT1_0 = "NO";
    defparam equal_152_0.INJECT1_1 = "YES";
    LUT4 i1_2_lut_3_lut_4_lut_adj_712 (.A(n2022[37]), .B(n2022[46]), .C(n4478[8]), 
         .D(n70862), .Z(n23081)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_712.init = 16'hf0e0;
    LUT4 i54366_3_lut (.A(\temp_outputs[2] [28]), .B(\temp_outputs[3] [28]), 
         .C(i[0]), .Z(n67277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54366_3_lut.init = 16'hcaca;
    LUT4 i54365_3_lut (.A(\temp_outputs[0] [28]), .B(\temp_outputs[1] [28]), 
         .C(i[0]), .Z(n67276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54365_3_lut.init = 16'hcaca;
    LUT4 i54363_3_lut (.A(\temp_outputs[2] [29]), .B(\temp_outputs[3] [29]), 
         .C(i[0]), .Z(n67274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54363_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_713 (.A(n2022[37]), .B(n2022[46]), .C(n4478[7]), 
         .D(n70862), .Z(n23090)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_713.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_714 (.A(n2022[37]), .B(n2022[46]), .C(n4478[6]), 
         .D(n70862), .Z(n23099)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_714.init = 16'hf0e0;
    CCU2D add_4584_add_1_add_1_13 (.A0(n14054), .B0(numL[0]), .C0(n12), 
          .D0(n921), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n61487), .S0(n3[11]));
    defparam add_4584_add_1_add_1_13.INIT0 = 16'hfe00;
    defparam add_4584_add_1_add_1_13.INIT1 = 16'h0000;
    defparam add_4584_add_1_add_1_13.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_715 (.A(n2022[37]), .B(n2022[46]), .C(n4478[5]), 
         .D(n70862), .Z(n23108)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_715.init = 16'hf0e0;
    LUT4 i54362_3_lut (.A(\temp_outputs[0] [29]), .B(\temp_outputs[1] [29]), 
         .C(i[0]), .Z(n67273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54362_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_716 (.A(n2022[37]), .B(n2022[46]), .C(n4478[4]), 
         .D(n70862), .Z(n23117)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_716.init = 16'hf0e0;
    LUT4 i54360_3_lut (.A(\temp_outputs[2] [30]), .B(\temp_outputs[3] [30]), 
         .C(i[0]), .Z(n67271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54360_3_lut.init = 16'hcaca;
    LUT4 i54359_3_lut (.A(\temp_outputs[0] [30]), .B(\temp_outputs[1] [30]), 
         .C(i[0]), .Z(n67270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54359_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_717 (.A(n2022[37]), .B(n2022[46]), .C(n4478[3]), 
         .D(n70862), .Z(n23126)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_717.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_718 (.A(n2022[37]), .B(n2022[46]), .C(n4478[2]), 
         .D(n70862), .Z(n22787)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_718.init = 16'hf0e0;
    LUT4 i54357_3_lut (.A(\temp_outputs[2] [31]), .B(\temp_outputs[3] [31]), 
         .C(i[0]), .Z(n67268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54357_3_lut.init = 16'hcaca;
    LUT4 i54356_3_lut (.A(\temp_outputs[0] [31]), .B(\temp_outputs[1] [31]), 
         .C(i[0]), .Z(n67267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54356_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_719 (.A(n2022[37]), .B(n2022[46]), .C(n4478[1]), 
         .D(n70862), .Z(n22796)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_719.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_720 (.A(n2022[37]), .B(n2022[46]), .C(n4478[26]), 
         .D(n70862), .Z(n23339)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_720.init = 16'hf0e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_721 (.A(n2022[37]), .B(n2022[46]), .C(n4478[24]), 
         .D(n70862), .Z(n23330)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_721.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_893 (.A(n2022[37]), .B(n2022[46]), .Z(n70863)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_893.init = 16'heeee;
    LUT4 i1_2_lut_rep_843_4_lut (.A(n2022[42]), .B(n2022[40]), .C(n2022[48]), 
         .D(n70863), .Z(n70813)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_843_4_lut.init = 16'hfffe;
    LUT4 i54354_3_lut (.A(\temp_outputs[2] [20]), .B(\temp_outputs[3] [20]), 
         .C(i[0]), .Z(n67265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54354_3_lut.init = 16'hcaca;
    LUT4 i54353_3_lut (.A(\temp_outputs[0] [20]), .B(\temp_outputs[1] [20]), 
         .C(i[0]), .Z(n67264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54353_3_lut.init = 16'hcaca;
    CCU2D add_4597_2 (.A0(i[0]), .B0(h[1]), .C0(GND_net), .D0(GND_net), 
          .A1(i[1]), .B1(h[2]), .C1(GND_net), .D1(GND_net), .COUT(n61477), 
          .S1(n7729[1]));
    defparam add_4597_2.INIT0 = 16'h7000;
    defparam add_4597_2.INIT1 = 16'h5666;
    defparam add_4597_2.INJECT1_0 = "NO";
    defparam add_4597_2.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_892 (.A(n2022[42]), .B(n2022[40]), .C(n2022[48]), 
         .Z(n70862)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_892.init = 16'hfefe;
    LUT4 i55006_2_lut (.A(o[0]), .B(\mlp_outputs[0] [31]), .Z(n67623)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i55006_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_722 (.A(\mlp_outputs[0] [31]), .B(n70809), .C(float_alu_c[31]), 
         .D(o[0]), .Z(n22859)) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_722.init = 16'h88c0;
    LUT4 i2_2_lut_rep_813_3_lut (.A(h[1]), .B(h[0]), .C(h[2]), .Z(n70783)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_rep_813_3_lut.init = 16'h1010;
    LUT4 i1_4_lut_adj_723 (.A(n32_adj_289), .B(n22859), .C(n2022[39]), 
         .D(n67623), .Z(n66434)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i1_4_lut_adj_723.init = 16'heefe;
    LUT4 i53911_2_lut_rep_891 (.A(h[1]), .B(h[0]), .Z(n70861)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i53911_2_lut_rep_891.init = 16'heeee;
    LUT4 i1_4_lut_adj_724 (.A(n11102[0]), .B(n61278[0]), .C(n2022[29]), 
         .D(n2022[7]), .Z(n6_adj_401)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_724.init = 16'heca0;
    LUT4 i1_2_lut_rep_890 (.A(n2022[13]), .B(n2022[35]), .Z(n70860)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_890.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_725 (.A(n2022[18]), .B(n2022[40]), .C(n70768), 
         .D(n70866), .Z(n23942)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_725.init = 16'h00fe;
    LUT4 i1_3_lut_4_lut_adj_726 (.A(n2022[18]), .B(n2022[40]), .C(n22276), 
         .D(n70866), .Z(n23975)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_726.init = 16'h00fe;
    CCU2D add_4597_4 (.A0(i[2]), .B0(h[3]), .C0(GND_net), .D0(GND_net), 
          .A1(\i[3] ), .B1(h[4]), .C1(GND_net), .D1(GND_net), .CIN(n61477), 
          .COUT(n61478), .S0(n7729[2]), .S1(n7729[3]));
    defparam add_4597_4.INIT0 = 16'h5666;
    defparam add_4597_4.INIT1 = 16'h5666;
    defparam add_4597_4.INJECT1_0 = "NO";
    defparam add_4597_4.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_889 (.A(n2022[18]), .B(n2022[40]), .Z(n70859)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_889.init = 16'heeee;
    LUT4 i2_2_lut_rep_755_3_lut_4_lut (.A(n2022[26]), .B(n2022[48]), .C(n70768), 
         .D(n22276), .Z(n70725)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_rep_755_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_727 (.A(n2022[26]), .B(n2022[48]), .C(n70866), 
         .D(n70860), .Z(n23977)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_727.init = 16'h0f0e;
    LUT4 i1_2_lut_3_lut_4_lut_adj_728 (.A(n2022[26]), .B(n2022[48]), .C(n2022[20]), 
         .D(n2022[42]), .Z(n22424)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_728.init = 16'hfffe;
    LUT4 i1_2_lut_rep_888 (.A(n2022[26]), .B(n2022[48]), .Z(n70858)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_888.init = 16'heeee;
    LUT4 i54348_3_lut (.A(\temp_outputs[2] [0]), .B(\temp_outputs[3] [0]), 
         .C(i[0]), .Z(n67259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54348_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_887 (.A(n2022[42]), .B(n2022[20]), .Z(n70857)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_887.init = 16'heeee;
    LUT4 i54347_3_lut (.A(\temp_outputs[0] [0]), .B(\temp_outputs[1] [0]), 
         .C(i[0]), .Z(n67258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54347_3_lut.init = 16'hcaca;
    LUT4 select_446_Select_0_i2_2_lut (.A(addr[0]), .B(n2022[1]), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam select_446_Select_0_i2_2_lut.init = 16'h8888;
    CCU2D equal_97_32 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n60978), 
          .S0(n1423));
    defparam equal_97_32.INIT0 = 16'hFFFF;
    defparam equal_97_32.INIT1 = 16'h0000;
    defparam equal_97_32.INJECT1_0 = "NO";
    defparam equal_97_32.INJECT1_1 = "NO";
    CCU2D add_4597_6 (.A0(\i[4] ), .B0(h[5]), .C0(GND_net), .D0(GND_net), 
          .A1(\i[5] ), .B1(h[6]), .C1(GND_net), .D1(GND_net), .CIN(n61478), 
          .COUT(n61479), .S0(n7729[4]), .S1(n7729[5]));
    defparam add_4597_6.INIT0 = 16'h5666;
    defparam add_4597_6.INIT1 = 16'h5666;
    defparam add_4597_6.INJECT1_0 = "NO";
    defparam add_4597_6.INJECT1_1 = "NO";
    CCU2D add_4597_8 (.A0(\i[6] ), .B0(h[7]), .C0(GND_net), .D0(GND_net), 
          .A1(\i[7] ), .B1(h[8]), .C1(GND_net), .D1(GND_net), .CIN(n61479), 
          .COUT(n61480), .S0(n7729[6]), .S1(n7729[7]));
    defparam add_4597_8.INIT0 = 16'h5666;
    defparam add_4597_8.INIT1 = 16'h5666;
    defparam add_4597_8.INJECT1_0 = "NO";
    defparam add_4597_8.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_729 (.A(mlp_done), .B(n3988), .C(n28181), 
         .Z(n66628)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_729.init = 16'h0808;
    LUT4 i2_3_lut_4_lut (.A(mlp_done), .B(n3988), .C(n28181), .D(SDA_c), 
         .Z(n23639)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0080;
    LUT4 i3_4_lut_adj_730 (.A(n3_adj_405[0]), .B(n6_adj_401), .C(n2022[32]), 
         .D(counter[0]), .Z(n8_adj_402)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B+(C (D)))) */ ;
    defparam i3_4_lut_adj_730.init = 16'hdcec;
    LUT4 i34472_1_lut_2_lut (.A(n2036), .B(mlp_mode), .Z(n3860)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i34472_1_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_878 (.A(n2036), .B(mlp_mode), .Z(n70848)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_878.init = 16'h2222;
    LUT4 i29987_2_lut_rep_821_3_lut (.A(h[2]), .B(h[1]), .C(h[0]), .Z(n70791)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i29987_2_lut_rep_821_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_819_3_lut (.A(h[2]), .B(h[1]), .C(h[0]), .Z(n70789)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_819_3_lut.init = 16'h1010;
    LUT4 i29418_2_lut_rep_877 (.A(h[2]), .B(h[1]), .Z(n70847)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i29418_2_lut_rep_877.init = 16'heeee;
    LUT4 i55105_3_lut_rep_725_3_lut_4_lut (.A(n2022[16]), .B(n2022[9]), 
         .C(n70822), .D(n70701), .Z(n70695)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i55105_3_lut_rep_725_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_rep_876 (.A(n2022[16]), .B(n2022[9]), .Z(n70846)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_876.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_731 (.A(\float_alu_mode[1] ), .B(\float_alu_mode[2] ), 
         .C(n1156), .D(n73809), .Z(n45598)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_731.init = 16'h8000;
    LUT4 i1_2_lut_rep_817_3_lut (.A(h[1]), .B(h[2]), .C(h[0]), .Z(n70787)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_rep_817_3_lut.init = 16'h0202;
    CCU2D add_4558_add_2_add_1_13 (.A0(o[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62765), .S0(n3_adj_405[11]));
    defparam add_4558_add_2_add_1_13.INIT0 = 16'hfaaa;
    defparam add_4558_add_2_add_1_13.INIT1 = 16'h0000;
    defparam add_4558_add_2_add_1_13.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_13.INJECT1_1 = "NO";
    CCU2D add_4558_add_2_add_1_11 (.A0(o[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62764), .COUT(n62765), .S0(n3_adj_405[9]), .S1(n3_adj_405[10]));
    defparam add_4558_add_2_add_1_11.INIT0 = 16'hfaaa;
    defparam add_4558_add_2_add_1_11.INIT1 = 16'hfaaa;
    defparam add_4558_add_2_add_1_11.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_11.INJECT1_1 = "NO";
    CCU2D add_4558_add_2_add_1_9 (.A0(o[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62763), .COUT(n62764), .S0(n3_adj_405[7]), .S1(n3_adj_405[8]));
    defparam add_4558_add_2_add_1_9.INIT0 = 16'hfaaa;
    defparam add_4558_add_2_add_1_9.INIT1 = 16'hfaaa;
    defparam add_4558_add_2_add_1_9.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_815_3_lut (.A(h[1]), .B(h[2]), .C(h[0]), .Z(n70785)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_815_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_875 (.A(h[1]), .B(h[2]), .Z(n70845)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_875.init = 16'h2222;
    CCU2D add_4558_add_2_add_1_7 (.A0(o[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62762), .COUT(n62763), .S0(n3_adj_405[5]), .S1(n3_adj_405[6]));
    defparam add_4558_add_2_add_1_7.INIT0 = 16'hfaaa;
    defparam add_4558_add_2_add_1_7.INIT1 = 16'hfaaa;
    defparam add_4558_add_2_add_1_7.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_7.INJECT1_1 = "NO";
    CCU2D add_4558_add_2_add_1_5 (.A0(o[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62761), .COUT(n62762), .S0(n3_adj_405[3]), .S1(n3_adj_405[4]));
    defparam add_4558_add_2_add_1_5.INIT0 = 16'hfaaa;
    defparam add_4558_add_2_add_1_5.INIT1 = 16'hfaaa;
    defparam add_4558_add_2_add_1_5.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_5.INJECT1_1 = "NO";
    CCU2D add_4558_add_2_add_1_3 (.A0(o[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62760), .COUT(n62761), .S0(n3_adj_405[1]), .S1(n3_adj_405[2]));
    defparam add_4558_add_2_add_1_3.INIT0 = 16'hfaaa;
    defparam add_4558_add_2_add_1_3.INIT1 = 16'h0555;
    defparam add_4558_add_2_add_1_3.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_3.INJECT1_1 = "NO";
    CCU2D add_4558_add_2_add_1_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n62760), .S1(n3_adj_405[0]));
    defparam add_4558_add_2_add_1_1.INIT0 = 16'hF000;
    defparam add_4558_add_2_add_1_1.INIT1 = 16'h0555;
    defparam add_4558_add_2_add_1_1.INJECT1_0 = "NO";
    defparam add_4558_add_2_add_1_1.INJECT1_1 = "NO";
    LUT4 i54345_3_lut (.A(\hidden_outputs[2] [0]), .B(\hidden_outputs[3] [0]), 
         .C(h[0]), .Z(n67256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54345_3_lut.init = 16'hcaca;
    LUT4 i54344_3_lut (.A(\hidden_outputs[0] [0]), .B(\hidden_outputs[1] [0]), 
         .C(h[0]), .Z(n67255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54344_3_lut.init = 16'hcaca;
    CCU2D add_4584_add_1_add_1_3 (.A0(n14054), .B0(numL[0]), .C0(n12), 
          .D0(n931), .A1(n13947[2]), .B1(n14054), .C1(numL[0]), .D1(n12), 
          .CIN(n61482), .COUT(n61483), .S0(n3[1]), .S1(n3[2]));
    defparam add_4584_add_1_add_1_3.INIT0 = 16'hfe00;
    defparam add_4584_add_1_add_1_3.INIT1 = 16'h5556;
    defparam add_4584_add_1_add_1_3.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_3.INJECT1_1 = "NO";
    CCU2D equal_97_32_49659 (.A0(\i[7] ), .B0(\i[6] ), .C0(\i[5] ), .D0(\i[4] ), 
          .A1(\i[4] ), .B1(\i[3] ), .C1(i[2]), .D1(i[1]), .CIN(n60977), 
          .COUT(n60978));
    defparam equal_97_32_49659.INIT0 = 16'h8001;
    defparam equal_97_32_49659.INIT1 = 16'h8001;
    defparam equal_97_32_49659.INJECT1_0 = "YES";
    defparam equal_97_32_49659.INJECT1_1 = "YES";
    LUT4 i4_4_lut_adj_732 (.A(n61250[0]), .B(n8_adj_402), .C(n2), .D(n2022[10]), 
         .Z(n63142)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i4_4_lut_adj_732.init = 16'hfefc;
    CCU2D add_4584_add_1_add_1_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n13947[0]), .B1(n14054), .C1(numL[0]), .D1(n12), 
          .COUT(n61482), .S1(n3[0]));
    defparam add_4584_add_1_add_1_1.INIT0 = 16'hF000;
    defparam add_4584_add_1_add_1_1.INIT1 = 16'h5556;
    defparam add_4584_add_1_add_1_1.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_733 (.A(n22276), .B(n23104), .C(n70862), .D(n70812), 
         .Z(n63026)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_733.init = 16'hfffe;
    LUT4 i1_3_lut_adj_734 (.A(n70866), .B(n63026), .C(float_alu_ready), 
         .Z(n27939)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i1_3_lut_adj_734.init = 16'heaea;
    LUT4 i54342_3_lut (.A(\hidden_outputs[2] [0]), .B(\hidden_outputs[3] [0]), 
         .C(n[0]), .Z(n67253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54342_3_lut.init = 16'hcaca;
    LUT4 i54341_3_lut (.A(\hidden_outputs[0] [0]), .B(\hidden_outputs[1] [0]), 
         .C(n[0]), .Z(n67252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i54341_3_lut.init = 16'hcaca;
    LUT4 i7119_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[9]), 
         .Z(n17905)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7119_2_lut_3_lut.init = 16'he0e0;
    LUT4 i49858_2_lut (.A(n3[0]), .B(h[0]), .Z(n61264[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49858_2_lut.init = 16'h6666;
    LUT4 i7117_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[10]), 
         .Z(n17901)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7117_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7112_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[13]), 
         .Z(n17891)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7112_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6918_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[14]), 
         .Z(n17567)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6918_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7110_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[15]), 
         .Z(n17887)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7110_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6685_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[16]), 
         .Z(n17309)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6685_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6717_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[17]), 
         .Z(n17345)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6717_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6735_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[18]), 
         .Z(n17365)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6735_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_33 (.A0(addr[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62711), .S0(n134_adj_408[31]));
    defparam addr_4653_add_4_33.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_33.INIT1 = 16'h0000;
    defparam addr_4653_add_4_33.INJECT1_0 = "NO";
    defparam addr_4653_add_4_33.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_31 (.A0(addr[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62710), .COUT(n62711), .S0(n134_adj_408[29]), .S1(n134_adj_408[30]));
    defparam addr_4653_add_4_31.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_31.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_31.INJECT1_0 = "NO";
    defparam addr_4653_add_4_31.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_29 (.A0(addr[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62709), .COUT(n62710), .S0(n134_adj_408[27]), .S1(n134_adj_408[28]));
    defparam addr_4653_add_4_29.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_29.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_29.INJECT1_0 = "NO";
    defparam addr_4653_add_4_29.INJECT1_1 = "NO";
    LUT4 i6771_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[19]), 
         .Z(n17405)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6771_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6952_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[20]), 
         .Z(n17619)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6952_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6963_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[21]), 
         .Z(n17634)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6963_2_lut_3_lut.init = 16'he0e0;
    LUT4 i53982_3_lut (.A(n70786), .B(numL[31]), .C(n66671), .Z(n66887)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i53982_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut_adj_735 (.A(n70723), .B(n4613), .C(numL[0]), .D(n66887), 
         .Z(n34857)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i3_4_lut_adj_735.init = 16'h0040;
    CCU2D addr_4653_add_4_27 (.A0(addr[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62708), .COUT(n62709), .S0(n134_adj_408[25]), .S1(n134_adj_408[26]));
    defparam addr_4653_add_4_27.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_27.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_27.INJECT1_0 = "NO";
    defparam addr_4653_add_4_27.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_25 (.A0(addr[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62707), .COUT(n62708), .S0(n134_adj_408[23]), .S1(n134_adj_408[24]));
    defparam addr_4653_add_4_25.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_25.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_25.INJECT1_0 = "NO";
    defparam addr_4653_add_4_25.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_23 (.A0(addr[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62706), .COUT(n62707), .S0(n134_adj_408[21]), .S1(n134_adj_408[22]));
    defparam addr_4653_add_4_23.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_23.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_23.INJECT1_0 = "NO";
    defparam addr_4653_add_4_23.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_21 (.A0(addr[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62705), .COUT(n62706), .S0(n134_adj_408[19]), .S1(n134_adj_408[20]));
    defparam addr_4653_add_4_21.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_21.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_21.INJECT1_0 = "NO";
    defparam addr_4653_add_4_21.INJECT1_1 = "NO";
    LUT4 i6965_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[22]), 
         .Z(n17638)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6965_2_lut_3_lut.init = 16'he0e0;
    LUT4 i6969_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[23]), 
         .Z(n17644)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6969_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7019_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[30]), 
         .Z(n17726)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7019_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7030_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n3998[31]), 
         .Z(n17745)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7030_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7528_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[0]), 
         .Z(n18717)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7528_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_19 (.A0(addr[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62704), .COUT(n62705), .S0(n134_adj_408[17]), .S1(n134_adj_408[18]));
    defparam addr_4653_add_4_19.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_19.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_19.INJECT1_0 = "NO";
    defparam addr_4653_add_4_19.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_17 (.A0(addr[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62703), .COUT(n62704), .S0(n134_adj_408[15]), .S1(n134_adj_408[16]));
    defparam addr_4653_add_4_17.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_17.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_17.INJECT1_0 = "NO";
    defparam addr_4653_add_4_17.INJECT1_1 = "NO";
    LUT4 i7005_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[28]), 
         .Z(n17704)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7005_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_15 (.A0(addr[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62702), .COUT(n62703), .S0(n134_adj_408[13]), .S1(n134_adj_408[14]));
    defparam addr_4653_add_4_15.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_15.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_15.INJECT1_0 = "NO";
    defparam addr_4653_add_4_15.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_13 (.A0(addr[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62701), .COUT(n62702), .S0(n134_adj_408[11]), .S1(n134_adj_408[12]));
    defparam addr_4653_add_4_13.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_13.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_13.INJECT1_0 = "NO";
    defparam addr_4653_add_4_13.INJECT1_1 = "NO";
    LUT4 i6972_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[24]), 
         .Z(n17650)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i6972_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7228_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[1]), 
         .Z(n18119)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7228_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7229_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[2]), 
         .Z(n18121)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7229_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_11 (.A0(addr[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62700), .COUT(n62701), .S0(n134_adj_408[9]), .S1(n134_adj_408[10]));
    defparam addr_4653_add_4_11.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_11.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_11.INJECT1_0 = "NO";
    defparam addr_4653_add_4_11.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_9 (.A0(addr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62699), .COUT(n62700), .S0(n134_adj_408[7]), .S1(n134_adj_408[8]));
    defparam addr_4653_add_4_9.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_9.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_9.INJECT1_0 = "NO";
    defparam addr_4653_add_4_9.INJECT1_1 = "NO";
    LUT4 i7129_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[3]), 
         .Z(n17925)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7129_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_7 (.A0(addr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62698), .COUT(n62699), .S0(n134_adj_408[5]), .S1(n134_adj_408[6]));
    defparam addr_4653_add_4_7.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_7.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_7.INJECT1_0 = "NO";
    defparam addr_4653_add_4_7.INJECT1_1 = "NO";
    CCU2D addr_4653_add_4_5 (.A0(addr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62697), .COUT(n62698), .S0(n134_adj_408[3]), .S1(n134_adj_408[4]));
    defparam addr_4653_add_4_5.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_5.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_5.INJECT1_0 = "NO";
    defparam addr_4653_add_4_5.INJECT1_1 = "NO";
    LUT4 i7127_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[4]), 
         .Z(n17921)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7127_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7126_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[5]), 
         .Z(n17919)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7126_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7107_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[6]), 
         .Z(n17881)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7107_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7122_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[7]), 
         .Z(n17911)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7122_2_lut_3_lut.init = 16'he0e0;
    LUT4 i7121_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[8]), 
         .Z(n17909)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7121_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_3 (.A0(addr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62696), .COUT(n62697), .S0(n134_adj_408[1]), .S1(n134_adj_408[2]));
    defparam addr_4653_add_4_3.INIT0 = 16'hfaaa;
    defparam addr_4653_add_4_3.INIT1 = 16'hfaaa;
    defparam addr_4653_add_4_3.INJECT1_0 = "NO";
    defparam addr_4653_add_4_3.INJECT1_1 = "NO";
    LUT4 i7116_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[11]), 
         .Z(n17899)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7116_2_lut_3_lut.init = 16'he0e0;
    CCU2D equal_97_30 (.A0(i_c[13]), .B0(\i[12] ), .C0(\i[11] ), .D0(i[10]), 
          .A1(i[10]), .B1(\i[9] ), .C1(\i[8] ), .D1(\i[7] ), .CIN(n60976), 
          .COUT(n60977));
    defparam equal_97_30.INIT0 = 16'h8001;
    defparam equal_97_30.INIT1 = 16'h8001;
    defparam equal_97_30.INJECT1_0 = "YES";
    defparam equal_97_30.INJECT1_1 = "YES";
    LUT4 i7114_2_lut_3_lut (.A(n2022[44]), .B(n2022[46]), .C(n4478[12]), 
         .Z(n17895)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7114_2_lut_3_lut.init = 16'he0e0;
    CCU2D addr_4653_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n62696), .S1(n134_adj_408[0]));
    defparam addr_4653_add_4_1.INIT0 = 16'hF000;
    defparam addr_4653_add_4_1.INIT1 = 16'h0555;
    defparam addr_4653_add_4_1.INJECT1_0 = "NO";
    defparam addr_4653_add_4_1.INJECT1_1 = "NO";
    LUT4 select_460_Select_0_i108_2_lut_rep_873 (.A(n2022[44]), .B(n2022[46]), 
         .Z(n70843)) /* synthesis lut_function=(A+(B)) */ ;
    defparam select_460_Select_0_i108_2_lut_rep_873.init = 16'heeee;
    CCU2D add_4584_add_1_add_1_9 (.A0(n14054), .B0(numL[0]), .C0(n12), 
          .D0(n925), .A1(n14054), .B1(numL[0]), .C1(n12), .D1(n924), 
          .CIN(n61485), .COUT(n61486), .S0(n3[7]), .S1(n3[8]));
    defparam add_4584_add_1_add_1_9.INIT0 = 16'hfe00;
    defparam add_4584_add_1_add_1_9.INIT1 = 16'hfe00;
    defparam add_4584_add_1_add_1_9.INJECT1_0 = "NO";
    defparam add_4584_add_1_add_1_9.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_32 (.A0(numL[30]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[31]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62694), .S0(n134_adj_407[30]), .S1(n134_adj_407[31]));
    defparam numL_4656_add_4_32.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_32.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_32.INJECT1_0 = "NO";
    defparam numL_4656_add_4_32.INJECT1_1 = "NO";
    LUT4 i29560_2_lut_3_lut (.A(n[0]), .B(n[1]), .C(\hidden_outputs[4] [27]), 
         .Z(n6_adj_249)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29560_2_lut_3_lut.init = 16'h1010;
    CCU2D numL_4656_add_4_30 (.A0(numL[28]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62693), .COUT(n62694), .S0(n134_adj_407[28]), .S1(n134_adj_407[29]));
    defparam numL_4656_add_4_30.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_30.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_30.INJECT1_0 = "NO";
    defparam numL_4656_add_4_30.INJECT1_1 = "NO";
    LUT4 i29562_2_lut_3_lut (.A(n[0]), .B(n[1]), .C(\hidden_outputs[4] [29]), 
         .Z(n6_adj_244)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29562_2_lut_3_lut.init = 16'h1010;
    CCU2D numL_4656_add_4_28 (.A0(numL[26]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62692), .COUT(n62693), .S0(n134_adj_407[26]), .S1(n134_adj_407[27]));
    defparam numL_4656_add_4_28.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_28.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_28.INJECT1_0 = "NO";
    defparam numL_4656_add_4_28.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_26 (.A0(numL[24]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62691), .COUT(n62692), .S0(n134_adj_407[24]), .S1(n134_adj_407[25]));
    defparam numL_4656_add_4_26.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_26.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_26.INJECT1_0 = "NO";
    defparam numL_4656_add_4_26.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_24 (.A0(numL[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62690), .COUT(n62691), .S0(n134_adj_407[22]), .S1(n134_adj_407[23]));
    defparam numL_4656_add_4_24.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_24.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_24.INJECT1_0 = "NO";
    defparam numL_4656_add_4_24.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_22 (.A0(numL[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62689), .COUT(n62690), .S0(n134_adj_407[20]), .S1(n134_adj_407[21]));
    defparam numL_4656_add_4_22.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_22.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_22.INJECT1_0 = "NO";
    defparam numL_4656_add_4_22.INJECT1_1 = "NO";
    LUT4 i29558_2_lut_3_lut (.A(n[0]), .B(n[1]), .C(\hidden_outputs[4] [25]), 
         .Z(n6_adj_259)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29558_2_lut_3_lut.init = 16'h1010;
    CCU2D numL_4656_add_4_20 (.A0(numL[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62688), .COUT(n62689), .S0(n134_adj_407[18]), .S1(n134_adj_407[19]));
    defparam numL_4656_add_4_20.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_20.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_20.INJECT1_0 = "NO";
    defparam numL_4656_add_4_20.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_18 (.A0(numL[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62687), .COUT(n62688), .S0(n134_adj_407[16]), .S1(n134_adj_407[17]));
    defparam numL_4656_add_4_18.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_18.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_18.INJECT1_0 = "NO";
    defparam numL_4656_add_4_18.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_16 (.A0(numL[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62686), .COUT(n62687), .S0(n134_adj_407[14]), .S1(n134_adj_407[15]));
    defparam numL_4656_add_4_16.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_16.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_16.INJECT1_0 = "NO";
    defparam numL_4656_add_4_16.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_14 (.A0(numL[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62685), .COUT(n62686), .S0(n134_adj_407[12]), .S1(n134_adj_407[13]));
    defparam numL_4656_add_4_14.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_14.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_14.INJECT1_0 = "NO";
    defparam numL_4656_add_4_14.INJECT1_1 = "NO";
    LUT4 i29559_2_lut_3_lut (.A(n[0]), .B(n[1]), .C(\hidden_outputs[4] [26]), 
         .Z(n6_adj_254)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i29559_2_lut_3_lut.init = 16'h1010;
    CCU2D numL_4656_add_4_12 (.A0(numL[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62684), .COUT(n62685), .S0(n134_adj_407[10]), .S1(n134_adj_407[11]));
    defparam numL_4656_add_4_12.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_12.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_12.INJECT1_0 = "NO";
    defparam numL_4656_add_4_12.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_10 (.A0(numL[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62683), .COUT(n62684), .S0(n134_adj_407[8]), .S1(n134_adj_407[9]));
    defparam numL_4656_add_4_10.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_10.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_10.INJECT1_0 = "NO";
    defparam numL_4656_add_4_10.INJECT1_1 = "NO";
    LUT4 i7052_2_lut_rep_872 (.A(n[0]), .B(n[1]), .Z(n70842)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7052_2_lut_rep_872.init = 16'heeee;
    CCU2D numL_4656_add_4_8 (.A0(numL[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62682), .COUT(n62683), .S0(n134_adj_407[6]), .S1(n134_adj_407[7]));
    defparam numL_4656_add_4_8.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_8.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_8.INJECT1_0 = "NO";
    defparam numL_4656_add_4_8.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_6 (.A0(numL[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62681), .COUT(n62682), .S0(n134_adj_407[4]), .S1(n134_adj_407[5]));
    defparam numL_4656_add_4_6.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_6.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_6.INJECT1_0 = "NO";
    defparam numL_4656_add_4_6.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_4 (.A0(numL[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(numL[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n62680), .COUT(n62681), .S0(n134_adj_407[2]), .S1(n134_adj_407[3]));
    defparam numL_4656_add_4_4.INIT0 = 16'hfaaa;
    defparam numL_4656_add_4_4.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_4.INJECT1_0 = "NO";
    defparam numL_4656_add_4_4.INJECT1_1 = "NO";
    CCU2D numL_4656_add_4_2 (.A0(n2664), .B0(numL[0]), .C0(GND_net), .D0(GND_net), 
          .A1(n14054), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n62680), 
          .S1(n134_adj_407[1]));
    defparam numL_4656_add_4_2.INIT0 = 16'h7000;
    defparam numL_4656_add_4_2.INIT1 = 16'hfaaa;
    defparam numL_4656_add_4_2.INJECT1_0 = "NO";
    defparam numL_4656_add_4_2.INJECT1_1 = "NO";
    CCU2D h_4657_add_4_33 (.A0(h[31]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n62678), 
          .S0(n134[31]));
    defparam h_4657_add_4_33.INIT0 = 16'hfaaa;
    defparam h_4657_add_4_33.INIT1 = 16'h0000;
    defparam h_4657_add_4_33.INJECT1_0 = "NO";
    defparam h_4657_add_4_33.INJECT1_1 = "NO";
    LUT4 mux_4578_i3_3_lut (.A(n7702[1]), .B(h[2]), .C(n70712), .Z(n13918[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_4578_i3_3_lut.init = 16'hcaca;
    LUT4 i49747_2_lut (.A(n236[1]), .B(n236[0]), .Z(n61391)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i49747_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module sram_dp
//

module sram_dp (sram_input_A, GND_net, sram_address_A, sram_address_B, 
            clock, sram_ready_A, sram_ready_B, VCC_net, SDA_c, sram_output_B);
    input [31:0]sram_input_A;
    input GND_net;
    input [11:0]sram_address_A;
    input [11:0]sram_address_B;
    input clock;
    input sram_ready_A;
    input sram_ready_B;
    input VCC_net;
    input SDA_c;
    output [31:0]sram_output_B;
    
    
    ram_dp_true ram_dq_true0 (.sram_input_A({sram_input_A}), .GND_net(GND_net), 
            .sram_address_A({sram_address_A}), .sram_address_B({sram_address_B}), 
            .clock(clock), .sram_ready_A(sram_ready_A), .sram_ready_B(sram_ready_B), 
            .VCC_net(VCC_net), .SDA_c(SDA_c), .sram_output_B({sram_output_B})) /* synthesis NGD_DRC_MASK=1 */ ;
    
endmodule
//
// Verilog Description of module ram_dp_true
//

module ram_dp_true (sram_input_A, GND_net, sram_address_A, sram_address_B, 
            clock, sram_ready_A, sram_ready_B, VCC_net, SDA_c, sram_output_B) /* synthesis NGD_DRC_MASK=1 */ ;
    input [31:0]sram_input_A;
    input GND_net;
    input [11:0]sram_address_A;
    input [11:0]sram_address_B;
    input clock;
    input sram_ready_A;
    input sram_ready_B;
    input VCC_net;
    input SDA_c;
    output [31:0]sram_output_B;
    
    
    DP8KC ram_dp_true_0_2_13 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[4]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[5]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[4]), .DOB1(sram_output_B[5])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_2_13.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_2_13.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_2_13.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_2_13.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_2_13.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_2_13.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_2_13.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_2_13.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_2_13.GSR = "ENABLED";
    defparam ram_dp_true_0_2_13.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_2_13.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_2_13.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_2_13.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_2_13.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_15_0 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[30]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[31]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[30]), .DOB1(sram_output_B[31])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_15_0.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_15_0.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_15_0.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_15_0.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_15_0.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_15_0.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_15_0.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_15_0.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_15_0.GSR = "ENABLED";
    defparam ram_dp_true_0_15_0.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_15_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_15_0.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_15_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_15_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_1_14 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[2]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[3]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[2]), .DOB1(sram_output_B[3])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_1_14.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_1_14.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_1_14.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_1_14.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_1_14.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_1_14.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_1_14.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_1_14.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_1_14.GSR = "ENABLED";
    defparam ram_dp_true_0_1_14.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_1_14.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_1_14.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_1_14.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_1_14.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_0_15 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[0]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[1]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[0]), .DOB1(sram_output_B[1])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_0_15.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_0_15.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_0_15.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_0_15.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_0_15.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_0_15.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_0_15.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_0_15.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_0_15.GSR = "ENABLED";
    defparam ram_dp_true_0_0_15.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_0_15.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_0_15.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_0_15.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_0_15.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_3_12 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[6]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[7]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[6]), .DOB1(sram_output_B[7])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_3_12.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_3_12.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_3_12.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_3_12.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_3_12.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_3_12.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_3_12.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_3_12.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_3_12.GSR = "ENABLED";
    defparam ram_dp_true_0_3_12.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_3_12.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_3_12.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_3_12.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_3_12.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_4_11 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[8]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[9]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[8]), .DOB1(sram_output_B[9])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_4_11.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_4_11.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_4_11.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_4_11.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_4_11.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_4_11.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_4_11.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_4_11.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_4_11.GSR = "ENABLED";
    defparam ram_dp_true_0_4_11.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_4_11.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_4_11.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_4_11.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_4_11.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_5_10 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[10]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[11]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[10]), .DOB1(sram_output_B[11])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_5_10.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_5_10.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_5_10.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_5_10.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_5_10.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_5_10.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_5_10.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_5_10.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_5_10.GSR = "ENABLED";
    defparam ram_dp_true_0_5_10.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_5_10.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_5_10.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_5_10.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_5_10.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_6_9 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[12]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[13]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[12]), .DOB1(sram_output_B[13])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_6_9.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_6_9.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_6_9.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_6_9.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_6_9.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_6_9.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_6_9.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_6_9.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_6_9.GSR = "ENABLED";
    defparam ram_dp_true_0_6_9.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_6_9.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_6_9.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_6_9.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_6_9.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_7_8 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[14]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[15]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[14]), .DOB1(sram_output_B[15])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_7_8.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_7_8.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_7_8.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_7_8.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_7_8.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_7_8.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_7_8.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_7_8.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_7_8.GSR = "ENABLED";
    defparam ram_dp_true_0_7_8.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_7_8.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_7_8.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_7_8.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_7_8.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_8_7 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[16]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[17]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[16]), .DOB1(sram_output_B[17])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_8_7.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_8_7.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_8_7.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_8_7.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_8_7.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_8_7.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_8_7.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_8_7.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_8_7.GSR = "ENABLED";
    defparam ram_dp_true_0_8_7.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_8_7.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_8_7.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_8_7.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_8_7.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_9_6 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[18]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[19]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[18]), .DOB1(sram_output_B[19])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_9_6.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_9_6.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_9_6.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_9_6.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_9_6.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_9_6.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_9_6.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_9_6.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_9_6.GSR = "ENABLED";
    defparam ram_dp_true_0_9_6.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_9_6.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_9_6.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_9_6.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_9_6.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_10_5 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[20]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[21]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[20]), .DOB1(sram_output_B[21])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_10_5.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_10_5.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_10_5.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_10_5.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_10_5.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_10_5.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_10_5.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_10_5.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_10_5.GSR = "ENABLED";
    defparam ram_dp_true_0_10_5.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_10_5.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_10_5.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_10_5.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_10_5.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_11_4 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[22]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[23]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[22]), .DOB1(sram_output_B[23])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_11_4.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_11_4.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_11_4.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_11_4.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_11_4.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_11_4.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_11_4.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_11_4.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_11_4.GSR = "ENABLED";
    defparam ram_dp_true_0_11_4.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_11_4.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_11_4.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_11_4.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_11_4.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_12_3 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[24]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[25]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[24]), .DOB1(sram_output_B[25])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_12_3.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_12_3.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_12_3.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_12_3.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_12_3.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_12_3.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_12_3.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_12_3.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_12_3.GSR = "ENABLED";
    defparam ram_dp_true_0_12_3.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_12_3.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_12_3.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_12_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_12_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_13_2 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[26]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[27]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[26]), .DOB1(sram_output_B[27])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_13_2.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_13_2.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_13_2.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_13_2.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_13_2.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_13_2.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_13_2.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_13_2.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_13_2.GSR = "ENABLED";
    defparam ram_dp_true_0_13_2.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_13_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_13_2.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_13_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_13_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC ram_dp_true_0_14_1 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(sram_input_A[28]), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(sram_input_A[29]), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(sram_address_A[0]), 
          .ADA2(sram_address_A[1]), .ADA3(sram_address_A[2]), .ADA4(sram_address_A[3]), 
          .ADA5(sram_address_A[4]), .ADA6(sram_address_A[5]), .ADA7(sram_address_A[6]), 
          .ADA8(sram_address_A[7]), .ADA9(sram_address_A[8]), .ADA10(sram_address_A[9]), 
          .ADA11(sram_address_A[10]), .ADA12(sram_address_A[11]), .CEA(sram_ready_A), 
          .OCEA(sram_ready_A), .CLKA(clock), .WEA(VCC_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(SDA_c), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(sram_address_B[0]), .ADB2(sram_address_B[1]), 
          .ADB3(sram_address_B[2]), .ADB4(sram_address_B[3]), .ADB5(sram_address_B[4]), 
          .ADB6(sram_address_B[5]), .ADB7(sram_address_B[6]), .ADB8(sram_address_B[7]), 
          .ADB9(sram_address_B[8]), .ADB10(sram_address_B[9]), .ADB11(sram_address_B[10]), 
          .ADB12(sram_address_B[11]), .CEB(sram_ready_B), .OCEB(sram_ready_B), 
          .CLKB(clock), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(SDA_c), .DOB0(sram_output_B[28]), .DOB1(sram_output_B[29])) /* synthesis MEM_LPC_FILE="ram_dp_true.lpc", MEM_INIT_FILE="INIT_ALL_0s", syn_instantiated=1 */ ;   // c:/users/yisong/documents/new/mlp/sram_dp_true.vhd(358[17:28])
    defparam ram_dp_true_0_14_1.DATA_WIDTH_A = 2;
    defparam ram_dp_true_0_14_1.DATA_WIDTH_B = 2;
    defparam ram_dp_true_0_14_1.REGMODE_A = "NOREG";
    defparam ram_dp_true_0_14_1.REGMODE_B = "NOREG";
    defparam ram_dp_true_0_14_1.CSDECODE_A = "0b000";
    defparam ram_dp_true_0_14_1.CSDECODE_B = "0b000";
    defparam ram_dp_true_0_14_1.WRITEMODE_A = "NORMAL";
    defparam ram_dp_true_0_14_1.WRITEMODE_B = "NORMAL";
    defparam ram_dp_true_0_14_1.GSR = "ENABLED";
    defparam ram_dp_true_0_14_1.RESETMODE = "ASYNC";
    defparam ram_dp_true_0_14_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam ram_dp_true_0_14_1.INIT_DATA = "STATIC";
    defparam ram_dp_true_0_14_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam ram_dp_true_0_14_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
